module encoder (b,c);
	output [0:0] c;

	input [0:0] b;

	reg [0:0] c;

	always @(b)
	begin
	end
endmodule
