module encoder (b,c);
	output [18:0] c;

	input [5:0] b;

	reg [18:0] c;

	always @(b)
	begin
		c[0] = b[0];
		c[1] = b[1];
		c[2] = b[2];
		c[3] = b[3];
		c[4] = b[4];
		c[5] = b[5];
		c[6] = b[0] ^ b[1] ^ b[4] ^ b[5];
		c[7] = b[4] ^ b[5];
		c[8] = b[2] ^ b[3] ^ b[5];
		c[9] = b[0] ^ b[3] ^ b[4];
		c[10] = b[1] ^ b[3] ^ b[4] ^ b[5];
		c[11] = b[2] ^ b[4];
		c[12] = b[0] ^ b[1] ^ b[5];
		c[13] = b[0] ^ b[1] ^ b[4] ^ b[5];
		c[14] = b[0] ^ b[3];
		c[15] = b[2] ^ b[4];
		c[16] = b[1] ^ b[3] ^ b[4];
		c[17] = b[1] ^ b[2] ^ b[4] ^ b[5];
		c[18] = b[1] ^ b[2] ^ b[3];
	end
endmodule
