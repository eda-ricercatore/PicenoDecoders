
module decoder ( cx, d );
  input [18:0] cx;
  output [5:0] d;
  wire   n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530;

  MUX2X1 U122 ( .B(n413), .A(n414), .S(cx[5]), .Y(d[5]) );
  NOR2X1 U123 ( .A(n415), .B(n416), .Y(n414) );
  MUX2X1 U124 ( .B(n417), .A(n418), .S(cx[4]), .Y(d[4]) );
  NOR2X1 U125 ( .A(n419), .B(n416), .Y(n418) );
  NAND2X1 U126 ( .A(n420), .B(n421), .Y(n416) );
  MUX2X1 U127 ( .B(n422), .A(n421), .S(n423), .Y(d[3]) );
  AND2X1 U128 ( .A(n420), .B(n424), .Y(n422) );
  INVX1 U129 ( .A(n425), .Y(n420) );
  NAND3X1 U130 ( .A(n426), .B(n427), .C(n428), .Y(n425) );
  MUX2X1 U131 ( .B(n429), .A(n430), .S(cx[2]), .Y(d[2]) );
  NOR2X1 U132 ( .A(n431), .B(n432), .Y(n430) );
  INVX1 U133 ( .A(n433), .Y(n429) );
  MUX2X1 U134 ( .B(n434), .A(n435), .S(n436), .Y(d[1]) );
  NOR2X1 U135 ( .A(n433), .B(n432), .Y(n434) );
  NAND2X1 U136 ( .A(n437), .B(n427), .Y(n432) );
  MUX2X1 U137 ( .B(n427), .A(n438), .S(cx[0]), .Y(d[0]) );
  AND2X1 U138 ( .A(n426), .B(n437), .Y(n438) );
  INVX1 U139 ( .A(n439), .Y(n437) );
  NAND3X1 U140 ( .A(n428), .B(n421), .C(n424), .Y(n439) );
  NOR2X1 U141 ( .A(n415), .B(n419), .Y(n424) );
  INVX1 U142 ( .A(n413), .Y(n419) );
  NAND3X1 U143 ( .A(n440), .B(n441), .C(n442), .Y(n413) );
  NOR2X1 U144 ( .A(n443), .B(n444), .Y(n442) );
  NAND2X1 U145 ( .A(n445), .B(n446), .Y(n444) );
  INVX1 U146 ( .A(n417), .Y(n415) );
  NAND3X1 U147 ( .A(n447), .B(n448), .C(n449), .Y(n417) );
  NOR2X1 U148 ( .A(n450), .B(n451), .Y(n449) );
  NAND2X1 U149 ( .A(n446), .B(n452), .Y(n451) );
  NAND3X1 U150 ( .A(n453), .B(n454), .C(n455), .Y(n450) );
  NOR2X1 U151 ( .A(n456), .B(n457), .Y(n448) );
  NOR2X1 U152 ( .A(n458), .B(n459), .Y(n447) );
  NAND3X1 U153 ( .A(n460), .B(n461), .C(n462), .Y(n421) );
  NOR2X1 U154 ( .A(n440), .B(n463), .Y(n462) );
  INVX1 U155 ( .A(n464), .Y(n428) );
  NAND3X1 U156 ( .A(n465), .B(n466), .C(n467), .Y(n464) );
  NOR2X1 U157 ( .A(n468), .B(n469), .Y(n467) );
  OAI21X1 U158 ( .A(n470), .B(n453), .C(n471), .Y(n469) );
  OAI21X1 U159 ( .A(n452), .B(n472), .C(n473), .Y(n471) );
  MUX2X1 U160 ( .B(n474), .A(n475), .S(n463), .Y(n472) );
  NAND2X1 U161 ( .A(n476), .B(n453), .Y(n474) );
  OAI21X1 U162 ( .A(n477), .B(n440), .C(n478), .Y(n468) );
  NAND2X1 U163 ( .A(n479), .B(n480), .Y(n478) );
  OAI21X1 U164 ( .A(n457), .B(n454), .C(n476), .Y(n480) );
  INVX1 U165 ( .A(n481), .Y(n477) );
  OAI22X1 U166 ( .A(n453), .B(n473), .C(n443), .D(n482), .Y(n481) );
  MUX2X1 U167 ( .B(n483), .A(n456), .S(n484), .Y(n466) );
  AND2X1 U168 ( .A(n485), .B(n486), .Y(n465) );
  MUX2X1 U169 ( .B(n487), .A(n470), .S(n457), .Y(n486) );
  NOR2X1 U170 ( .A(n452), .B(n456), .Y(n487) );
  MUX2X1 U171 ( .B(n488), .A(n489), .S(n490), .Y(n485) );
  NAND2X1 U172 ( .A(n491), .B(n492), .Y(n489) );
  AOI22X1 U173 ( .A(n445), .B(n493), .C(n455), .D(n453), .Y(n492) );
  AOI22X1 U174 ( .A(n482), .B(n475), .C(n440), .D(n494), .Y(n491) );
  OAI21X1 U175 ( .A(n473), .B(n479), .C(n495), .Y(n488) );
  INVX1 U176 ( .A(n459), .Y(n495) );
  NAND3X1 U177 ( .A(n494), .B(n470), .C(n475), .Y(n459) );
  NOR2X1 U178 ( .A(n431), .B(n433), .Y(n426) );
  NOR2X1 U179 ( .A(n496), .B(n497), .Y(n433) );
  NAND3X1 U180 ( .A(n463), .B(n440), .C(n498), .Y(n497) );
  NAND3X1 U181 ( .A(n490), .B(n461), .C(n499), .Y(n496) );
  NOR2X1 U182 ( .A(n473), .B(n500), .Y(n499) );
  INVX1 U183 ( .A(n501), .Y(n461) );
  NAND3X1 U184 ( .A(n484), .B(n483), .C(n502), .Y(n501) );
  NOR2X1 U185 ( .A(n456), .B(n503), .Y(n502) );
  NAND2X1 U186 ( .A(n443), .B(n445), .Y(n503) );
  INVX1 U187 ( .A(n435), .Y(n431) );
  NAND3X1 U188 ( .A(n490), .B(n441), .C(n504), .Y(n435) );
  NOR2X1 U189 ( .A(n445), .B(n505), .Y(n504) );
  NAND2X1 U190 ( .A(n443), .B(n454), .Y(n505) );
  NOR2X1 U191 ( .A(n506), .B(n507), .Y(n441) );
  NAND3X1 U192 ( .A(n500), .B(n473), .C(n498), .Y(n507) );
  NOR3X1 U193 ( .A(n457), .B(n508), .C(n453), .Y(n498) );
  NAND3X1 U194 ( .A(n456), .B(n494), .C(n509), .Y(n506) );
  NOR2X1 U195 ( .A(n483), .B(n484), .Y(n509) );
  INVX1 U196 ( .A(n476), .Y(n484) );
  INVX1 U197 ( .A(n493), .Y(n483) );
  OR2X1 U198 ( .A(n510), .B(n511), .Y(n427) );
  NAND3X1 U199 ( .A(n463), .B(n460), .C(n440), .Y(n511) );
  INVX1 U200 ( .A(n454), .Y(n440) );
  XOR2X1 U201 ( .A(n512), .B(n513), .Y(n454) );
  XOR2X1 U202 ( .A(cx[8]), .B(cx[5]), .Y(n513) );
  NOR2X1 U203 ( .A(n514), .B(n515), .Y(n460) );
  NAND3X1 U204 ( .A(n500), .B(n473), .C(n508), .Y(n515) );
  INVX1 U205 ( .A(n470), .Y(n508) );
  XOR2X1 U206 ( .A(cx[4]), .B(n516), .Y(n470) );
  XOR2X1 U207 ( .A(cx[7]), .B(cx[5]), .Y(n516) );
  INVX1 U208 ( .A(n455), .Y(n473) );
  XNOR2X1 U209 ( .A(n517), .B(cx[13]), .Y(n455) );
  INVX1 U210 ( .A(n452), .Y(n500) );
  XNOR2X1 U211 ( .A(n518), .B(n519), .Y(n452) );
  XNOR2X1 U212 ( .A(cx[4]), .B(cx[9]), .Y(n518) );
  NAND3X1 U213 ( .A(n453), .B(n457), .C(n490), .Y(n514) );
  INVX1 U214 ( .A(n446), .Y(n490) );
  XNOR2X1 U215 ( .A(n520), .B(n521), .Y(n446) );
  XOR2X1 U216 ( .A(cx[17]), .B(n522), .Y(n521) );
  XNOR2X1 U217 ( .A(cx[2]), .B(cx[5]), .Y(n520) );
  XNOR2X1 U218 ( .A(n523), .B(n524), .Y(n457) );
  XOR2X1 U219 ( .A(cx[5]), .B(cx[10]), .Y(n524) );
  XNOR2X1 U220 ( .A(n525), .B(cx[15]), .Y(n453) );
  INVX1 U221 ( .A(n494), .Y(n463) );
  XOR2X1 U222 ( .A(n519), .B(cx[14]), .Y(n494) );
  XNOR2X1 U223 ( .A(cx[0]), .B(n423), .Y(n519) );
  NAND3X1 U224 ( .A(n475), .B(n456), .C(n526), .Y(n510) );
  INVX1 U225 ( .A(n458), .Y(n526) );
  NAND3X1 U226 ( .A(n476), .B(n493), .C(n479), .Y(n458) );
  INVX1 U227 ( .A(n445), .Y(n479) );
  XNOR2X1 U228 ( .A(n523), .B(cx[16]), .Y(n445) );
  XNOR2X1 U229 ( .A(cx[3]), .B(n522), .Y(n523) );
  XNOR2X1 U230 ( .A(n525), .B(cx[11]), .Y(n493) );
  XNOR2X1 U231 ( .A(cx[2]), .B(cx[4]), .Y(n525) );
  XNOR2X1 U232 ( .A(n527), .B(n512), .Y(n476) );
  XNOR2X1 U233 ( .A(cx[2]), .B(n423), .Y(n512) );
  INVX1 U234 ( .A(cx[3]), .Y(n423) );
  XNOR2X1 U235 ( .A(cx[1]), .B(cx[18]), .Y(n527) );
  INVX1 U236 ( .A(n482), .Y(n456) );
  XOR2X1 U237 ( .A(n528), .B(n529), .Y(n482) );
  XNOR2X1 U238 ( .A(cx[5]), .B(n436), .Y(n529) );
  XNOR2X1 U239 ( .A(cx[0]), .B(cx[12]), .Y(n528) );
  INVX1 U240 ( .A(n443), .Y(n475) );
  XNOR2X1 U241 ( .A(n517), .B(cx[6]), .Y(n443) );
  XOR2X1 U242 ( .A(n530), .B(n522), .Y(n517) );
  XNOR2X1 U243 ( .A(n436), .B(cx[4]), .Y(n522) );
  INVX1 U244 ( .A(cx[1]), .Y(n436) );
  XNOR2X1 U245 ( .A(cx[0]), .B(cx[5]), .Y(n530) );
endmodule

