`timescale 1ns/100ps
/**
 * `timescale time_unit base / precision base
 *
 * -Specifies the time units and precision for delays:
 * -time_unit is the amount of time a delay of 1 represents.
 *	The time unit must be 1 10 or 100
 * -base is the time base for each unit, ranging from seconds
 *	to femtoseconds, and must be: s ms us ns ps or fs
 * -precision and base represent how many decimal points of
 *	precision to use relative to the time units.
 */

/**
 * This is written by Zhiyang Ong -student number 6004919412-
 * for EE577b Homework 2, Question 2
 */

// Testbench for behavioral model for the decoder


// Import the modules that will be tested for in this testbench
`include "decoder4to16.v"

// IMPORTANT: To run this, try: ncverilog -f ee577bHw2q2.f +gui
module tb_decoder4to16();
	/**
	 * Declare signal types for testbench to drive and monitor
	 * signals during the simulation of the arbiter
	 *
	 * The reg data type holds a value until a new value is driven
	 * onto it in an "initial" or "always" block. It can only be
	 * assigned a value in an "always" or "initial" block, and is
	 * used to apply stimulus to the inputs of the DUT.
	 *
	 * The wire type is a passive data type that holds a value driven
	 * onto it by a port, assign statement or reg type. Wires cannot be
	 * assigned values inside "always" and "initial" blocks. They can
	 * be used to hold the values of the DUT's outputs
	 */
	
	// Declare "wire" signals: outputs from the DUT
	wire [15:1] dout;
	
	// Declare "reg" signals: inputs to the DUT
	reg [3:0] din;
	
	
	
	/**
	 * Instantiate an instance of arbiter_LRU4 so that
	 * inputs can be passed to the Device Under Test (DUT)
	 * Given instance name is "arb"
	 */
	decoder4to16 dec4to16 (
		// instance_name(signal name),
		// Signal name can be the same as the instance name
		din,dout);
	

	
	/**
	 * Initial block start executing sequentially @ t=0
	 * If and when a delay is encountered, the execution of this block
	 * pauses or waits until the delay time has passed, before resuming
	 * execution
	 *
	 * Each intial or always block executes concurrently; that is,
	 * multiple "always" or "initial" blocks will execute simultaneously
	 *
	 * E.g.
	 * always
	 * begin
	 *		#10 clk_50 = ~clk_50; // Invert clock signal every 10 ns
	 *		// Clock signal has a period of 20 ns or 50 MHz
	 * end
	 */
	initial
	begin
		// "$time" indicates the current time in the simulation
		$display(" << Starting the simulation >>");
		din = 15'd0;
		#1;
		din = 15'd1;
		
		// @ t=0,
		#1;
		din = 15'd2;
		
		
		#1;
		din = 15'd3;
		
				
		#1;
		din = 15'd4;
		
		#1;
		din = 15'd5;
		
		#1;
		din = 15'd6;
		
		#1;
		din = 15'd7;
		
		#1;
		din = 15'd8;
		
		#1;
		din = 15'd9;
		
		#1;
		din = 15'd10;

		#1;
		din = 15'd11;

		#1;
		din = 15'd12;

		#1;
		din = 15'd13;

		#1;
		din = 15'd14;

		#1;
		din = 15'd15;

		
		
				
		#20;
		
		$display(" << Finishing the simulation >>");
		$finish;
	end

endmodule
