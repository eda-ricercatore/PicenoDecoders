* # FILE NAME: /HOME/SCF-07/ZHIYANGO/SIMULATION/VITERBI_DECODER/HSPICES/        
* SCHEMATIC/NETLIST/VITERBI_DECODER.C.RAW
* NETLIST OUTPUT FOR HSPICES.
* GENERATED ON NOV 7 08:54:31 2007
   
* GLOBAL NET DEFINITIONS
.GLOBAL VDD! GND! VDD! 
* FILE NAME: VITERBI_VITERBI_DECODER_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: VITERBI_DECODER.
* GENERATED FOR: HSPICES.
* GENERATED ON NOV  7 08:54:36 2007.
   
XACS3 BRCH_MET5_1 BRCH_MET5_0 BRCH_MET7_1 BRCH_MET7_0 D3 N_PM3_3 N_PM3_2 
+N_PM3_1 N_PM3_0 P_M2_3 P_M2_2 P_M2_1 P_M2_0 P_M3_3 P_M3_2 P_M3_1 P_M3_0 SUB1 
XACS1 BRCH_MET4_1 BRCH_MET4_0 BRCH_MET6_1 BRCH_MET6_0 D1 N_PM1_3 N_PM1_2 
+N_PM1_1 N_PM1_0 P_M2_3 P_M2_2 P_M2_1 P_M2_0 P_M3_3 P_M3_2 P_M3_1 P_M3_0 SUB2 
XACS2 BRCH_MET1_1 BRCH_MET1_0 BRCH_MET3_1 BRCH_MET3_0 D2 N_PM2_3 N_PM2_2 
+N_PM2_1 N_PM2_0 P_M0_3 P_M0_2 P_M0_1 P_M0_0 P_M1_3 P_M1_2 P_M1_1 P_M1_0 SUB3 
XACS0 BRCH_MET0_1 BRCH_MET0_0 BRCH_MET2_1 BRCH_MET2_0 D0 N_PM0_3 N_PM0_2 
+N_PM0_1 N_PM0_0 P_M0_3 P_M0_2 P_M0_1 P_M0_0 P_M1_3 P_M1_2 P_M1_1 P_M1_0 SUB4 
XPATH_METRIC_SM CLK N_PM0_3 N_PM0_2 N_PM0_1 N_PM0_0 N_PM1_3 N_PM1_2 N_PM1_1 
+N_PM1_0 N_PM2_3 N_PM2_2 N_PM2_1 N_PM2_0 N_PM3_3 N_PM3_2 N_PM3_1 N_PM3_0 P_M0_3 
+P_M0_2 P_M0_1 P_M0_0 P_M1_3 P_M1_2 P_M1_1 P_M1_0 P_M2_3 P_M2_2 P_M2_1 P_M2_0 
+P_M3_3 P_M3_2 P_M3_1 P_M3_0 RESET PMSM_G32 
X0 CLK D0 D1 D2 D3 D P_M0_3 P_M0_2 P_M0_1 P_M0_0 P_M1_3 P_M1_2 P_M1_1 P_M1_0 
+P_M2_3 P_M2_2 P_M2_1 P_M2_0 P_M3_3 P_M3_2 P_M3_1 P_M3_0 RESET SPD_G33 
XBRCH_MET BRCH_MET0_1 BRCH_MET0_0 BRCH_MET1_1 BRCH_MET1_0 BRCH_MET2_1 
+BRCH_MET2_0 BRCH_MET3_1 BRCH_MET3_0 BRCH_MET4_1 BRCH_MET4_0 BRCH_MET5_1 
+BRCH_MET5_0 BRCH_MET6_1 BRCH_MET6_0 BRCH_MET7_1 BRCH_MET7_0 CX_0 CX_1 BMU_G34 
   
   
   
   
* FILE NAME: VITERBI_SPDU_2_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: SPDU_2.
* GENERATED FOR: HSPICES.
* GENERATED ON NOV  7 08:54:34 2007.
   
* TERMINAL MAPPING: CLK = CLK
*                   D0 = D0
*                   D1 = D1
*                   D2 = D2
*                   D3 = D3
*                   IN0 = IN0
*                   IN1 = IN1
*                   IN2 = IN2
*                   IN3 = IN3
*                   OUT0 = OUT0
*                   OUT1 = OUT1
*                   OUT2 = OUT2
*                   OUT3 = OUT3
*                   RESET = RESET
.SUBCKT SPDU_2_G18 CLK D0 D1 D2 D3 IN0 IN1 IN2 IN3 OUT0 OUT1 OUT2 OUT3 RESET 
XOUT1_REG CLK OUT1211 OUT1 DFFPOSX1_G14 
XOUT0_REG CLK OUT0205 OUT0 DFFPOSX1_G14 
XOUT2_REG CLK OUT2217 OUT2 DFFPOSX1_G14 
XOUT3_REG CLK OUT3223 OUT3 DFFPOSX1_G14 
XU37 RESET N1 OUT3223 NOR2X1_G7 
XU43 RESET N4 OUT0205 NOR2X1_G7 
XU41 RESET N3 OUT1211 NOR2X1_G7 
XU39 RESET N2 OUT2217 NOR2X1_G7 
XU38 IN3 IN2 D3 N1 MUX2X1_G5 
XU40 IN1 IN0 D2 N2 MUX2X1_G5 
XU42 IN3 IN2 D1 N3 MUX2X1_G5 
XU44 IN1 IN0 D0 N4 MUX2X1_G5 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS SPDU_2_G18 
* FILE NAME: VITERBI_SPDU_12_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: SPDU_12.
* GENERATED FOR: HSPICES.
* GENERATED ON NOV  7 08:54:35 2007.
   
* TERMINAL MAPPING: CLK = CLK
*                   D0 = D0
*                   D1 = D1
*                   D2 = D2
*                   D3 = D3
*                   IN0 = IN0
*                   IN1 = IN1
*                   IN2 = IN2
*                   IN3 = IN3
*                   OUT0 = OUT0
*                   OUT1 = OUT1
*                   OUT2 = OUT2
*                   OUT3 = OUT3
*                   RESET = RESET
.SUBCKT SPDU_12_G28 CLK D0 D1 D2 D3 IN0 IN1 IN2 IN3 OUT0 OUT1 OUT2 OUT3 RESET 
XOUT1_REG CLK OUT1211 OUT1 DFFPOSX1_G14 
XOUT2_REG CLK OUT2217 OUT2 DFFPOSX1_G14 
XOUT0_REG CLK OUT0205 OUT0 DFFPOSX1_G14 
XOUT3_REG CLK OUT3223 OUT3 DFFPOSX1_G14 
XU43 RESET N4 OUT0205 NOR2X1_G7 
XU39 RESET N2 OUT2217 NOR2X1_G7 
XU41 RESET N3 OUT1211 NOR2X1_G7 
XU37 RESET N1 OUT3223 NOR2X1_G7 
XU38 IN3 IN2 D3 N1 MUX2X1_G5 
XU40 IN1 IN0 D2 N2 MUX2X1_G5 
XU42 IN3 IN2 D1 N3 MUX2X1_G5 
XU44 IN1 IN0 D0 N4 MUX2X1_G5 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS SPDU_12_G28 
* FILE NAME: VITERBI_SPDU_5_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: SPDU_5.
* GENERATED FOR: HSPICES.
* GENERATED ON NOV  7 08:54:35 2007.
   
* TERMINAL MAPPING: CLK = CLK
*                   D0 = D0
*                   D1 = D1
*                   D2 = D2
*                   D3 = D3
*                   IN0 = IN0
*                   IN1 = IN1
*                   IN2 = IN2
*                   IN3 = IN3
*                   OUT0 = OUT0
*                   OUT1 = OUT1
*                   OUT2 = OUT2
*                   OUT3 = OUT3
*                   RESET = RESET
.SUBCKT SPDU_5_G26 CLK D0 D1 D2 D3 IN0 IN1 IN2 IN3 OUT0 OUT1 OUT2 OUT3 RESET 
XOUT2_REG CLK OUT2217 OUT2 DFFPOSX1_G14 
XOUT1_REG CLK OUT1211 OUT1 DFFPOSX1_G14 
XOUT3_REG CLK OUT3223 OUT3 DFFPOSX1_G14 
XOUT0_REG CLK OUT0205 OUT0 DFFPOSX1_G14 
XU37 RESET N1 OUT3223 NOR2X1_G7 
XU43 RESET N4 OUT0205 NOR2X1_G7 
XU39 RESET N2 OUT2217 NOR2X1_G7 
XU41 RESET N3 OUT1211 NOR2X1_G7 
XU38 IN3 IN2 D3 N1 MUX2X1_G5 
XU40 IN1 IN0 D2 N2 MUX2X1_G5 
XU44 IN1 IN0 D0 N4 MUX2X1_G5 
XU42 IN3 IN2 D1 N3 MUX2X1_G5 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS SPDU_5_G26 
* FILE NAME: OSU_STDCELLS_AND2X1_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: AND2X1.
* GENERATED FOR: HSPICES.
* GENERATED ON NOV  7 08:54:32 2007.
   
* TERMINAL MAPPING: A = A
*                   B = B
*                   Y = Y
.SUBCKT AND2X1_G8 A B Y 
M13 NET12 A VDD! VDD!  TSMC20P  L=200E-9 W=2E-6 AD=1E-12 AS=1E-12 PD=5E-6 
+PS=5E-6 M=1 
M14 NET12 B VDD! VDD!  TSMC20P  L=200E-9 W=2E-6 AD=1E-12 AS=1E-12 PD=5E-6 
+PS=5E-6 M=1 
M15 Y NET12 VDD! VDD!  TSMC20P  L=200E-9 W=2E-6 AD=1E-12 AS=1E-12 PD=5E-6 
+PS=5E-6 M=1 
M16 NET12 A NET15 0  TSMC20N  L=200E-9 W=2E-6 AD=1E-12 AS=1E-12 PD=5E-6 
+PS=5E-6 M=1 
M17 NET15 B 0 0  TSMC20N  L=200E-9 W=2E-6 AD=1E-12 AS=1E-12 PD=5E-6 PS=5E-6 
+M=1 
M18 Y NET12 0 0  TSMC20N  L=200E-9 W=1E-6 AD=500E-15 AS=500E-15 PD=3E-6 
+PS=3E-6 M=1 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS AND2X1_G8 
* FILE NAME: OSU_STDCELLS_NAND3X1_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: NAND3X1.
* GENERATED FOR: HSPICES.
* GENERATED ON NOV  7 08:54:33 2007.
   
* TERMINAL MAPPING: A = A
*                   B = B
*                   C = C
*                   Y = Y
.SUBCKT NAND3X1_G11 A B C Y 
M14 Y A NET9 0  TSMC20N  L=200E-9 W=3E-6 AD=1.5E-12 AS=1.5E-12 PD=7E-6 PS=7E-6 
+M=1 
M17 NET9 B NET013 0  TSMC20N  L=200E-9 W=3E-6 AD=1.5E-12 AS=1.5E-12 PD=7E-6 
+PS=7E-6 M=1 
M18 NET013 C 0 0  TSMC20N  L=200E-9 W=3E-6 AD=1.5E-12 AS=1.5E-12 PD=7E-6 
+PS=7E-6 M=1 
M13 Y A VDD! VDD!  TSMC20P  L=200E-9 W=2E-6 AD=1E-12 AS=1E-12 PD=5E-6 PS=5E-6 
+M=1 
M15 Y B VDD! VDD!  TSMC20P  L=200E-9 W=2E-6 AD=1E-12 AS=1E-12 PD=5E-6 PS=5E-6 
+M=1 
M16 Y C VDD! VDD!  TSMC20P  L=200E-9 W=2E-6 AD=1E-12 AS=1E-12 PD=5E-6 PS=5E-6 
+M=1 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS NAND3X1_G11 
* FILE NAME: VITERBI_SPDU_6_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: SPDU_6.
* GENERATED FOR: HSPICES.
* GENERATED ON NOV  7 08:54:34 2007.
   
* TERMINAL MAPPING: CLK = CLK
*                   D0 = D0
*                   D1 = D1
*                   D2 = D2
*                   D3 = D3
*                   IN0 = IN0
*                   IN1 = IN1
*                   IN2 = IN2
*                   IN3 = IN3
*                   OUT0 = OUT0
*                   OUT1 = OUT1
*                   OUT2 = OUT2
*                   OUT3 = OUT3
*                   RESET = RESET
.SUBCKT SPDU_6_G22 CLK D0 D1 D2 D3 IN0 IN1 IN2 IN3 OUT0 OUT1 OUT2 OUT3 RESET 
XOUT1_REG CLK OUT1211 OUT1 DFFPOSX1_G14 
XOUT3_REG CLK OUT3223 OUT3 DFFPOSX1_G14 
XOUT2_REG CLK OUT2217 OUT2 DFFPOSX1_G14 
XOUT0_REG CLK OUT0205 OUT0 DFFPOSX1_G14 
XU39 RESET N2 OUT2217 NOR2X1_G7 
XU41 RESET N3 OUT1211 NOR2X1_G7 
XU37 RESET N1 OUT3223 NOR2X1_G7 
XU43 RESET N4 OUT0205 NOR2X1_G7 
XU38 IN3 IN2 D3 N1 MUX2X1_G5 
XU44 IN1 IN0 D0 N4 MUX2X1_G5 
XU40 IN1 IN0 D2 N2 MUX2X1_G5 
XU42 IN3 IN2 D1 N3 MUX2X1_G5 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS SPDU_6_G22 
* FILE NAME: OSU_STDCELLS_LATCH_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: LATCH.
* GENERATED FOR: HSPICES.
* GENERATED ON NOV  7 08:54:33 2007.
   
* TERMINAL MAPPING: CLK = CLK
*                   D = D
*                   Q = Q
.SUBCKT LATCH_G12 CLK D Q 
M36 NET9 Q 0 0  TSMC20N  L=200E-9 W=1E-6 AD=500E-15 AS=500E-15 PD=3E-6 PS=3E-6 
+M=1 
M33 NET18 NET21 NET9 0  TSMC20N  L=200E-9 W=1E-6 AD=500E-15 AS=500E-15 PD=3E-6 
+PS=3E-6 M=1 
M32 NET18 CLK NET15 0  TSMC20N  L=200E-9 W=1E-6 AD=500E-15 AS=500E-15 PD=3E-6 
+PS=3E-6 M=1 
M35 Q NET18 0 0  TSMC20N  L=200E-9 W=2E-6 AD=1E-12 AS=1E-12 PD=5E-6 PS=5E-6 
+M=1 
M31 NET21 CLK 0 0  TSMC20N  L=200E-9 W=2E-6 AD=1E-12 AS=1E-12 PD=5E-6 PS=5E-6 
+M=1 
M34 NET15 D 0 0  TSMC20N  L=200E-9 W=1E-6 AD=500E-15 AS=500E-15 PD=3E-6 
+PS=3E-6 M=1 
M21 NET21 CLK VDD! VDD!  TSMC20P  L=200E-9 W=4E-6 AD=2E-12 AS=2E-12 PD=9E-6 
+PS=9E-6 M=1 
M26 NET35 Q VDD! VDD!  TSMC20P  L=200E-9 W=1E-6 AD=500E-15 AS=500E-15 PD=3E-6 
+PS=3E-6 M=1 
M27 NET26 D VDD! VDD!  TSMC20P  L=200E-9 W=2E-6 AD=1E-12 AS=1E-12 PD=5E-6 
+PS=5E-6 M=1 
M28 Q NET18 VDD! VDD!  TSMC20P  L=200E-9 W=4E-6 AD=2E-12 AS=2E-12 PD=9E-6 
+PS=9E-6 M=1 
M29 NET18 CLK NET35 VDD!  TSMC20P  L=200E-9 W=1E-6 AD=500E-15 AS=500E-15 
+PD=3E-6 PS=3E-6 M=1 
M30 NET18 NET21 NET26 VDD!  TSMC20P  L=200E-9 W=2E-6 AD=1E-12 AS=1E-12 PD=5E-6 
+PS=5E-6 M=1 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS LATCH_G12 
* FILE NAME: VITERBI_DEMUX_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: DEMUX.
* GENERATED FOR: HSPICES.
* GENERATED ON NOV  7 08:54:34 2007.
   
* TERMINAL MAPPING: D0 = D0
*                   D1 = D1
*                   IN0 = IN0
*                   IN1 = IN1
*                   IN2 = IN2
*                   IN3 = IN3
*                   OUT = OUT
.SUBCKT DEMUX_G15 D0 D1 IN0 IN1 IN2 IN3 OUT 
XU26 N2 N1 D1 OUT MUX2X1_G5 
XU27 IN3 IN2 D0 N2 MUX2X1_G5 
XU28 IN1 IN0 D0 N1 MUX2X1_G5 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS DEMUX_G15 
* FILE NAME: VITERBI_PMSM_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: PMSM.
* GENERATED FOR: HSPICES.
* GENERATED ON NOV  7 08:54:33 2007.
   
* TERMINAL MAPPING: CLK = CLK
*                   NPM0<3> = NPM0_3
*                   NPM0<2> = NPM0_2
*                   NPM0<1> = NPM0_1
*                   NPM0<0> = NPM0_0
*                   NPM1<3> = NPM1_3
*                   NPM1<2> = NPM1_2
*                   NPM1<1> = NPM1_1
*                   NPM1<0> = NPM1_0
*                   NPM2<3> = NPM2_3
*                   NPM2<2> = NPM2_2
*                   NPM2<1> = NPM2_1
*                   NPM2<0> = NPM2_0
*                   NPM3<3> = NPM3_3
*                   NPM3<2> = NPM3_2
*                   NPM3<1> = NPM3_1
*                   NPM3<0> = NPM3_0
*                   PM0<3> = PM0_3
*                   PM0<2> = PM0_2
*                   PM0<1> = PM0_1
*                   PM0<0> = PM0_0
*                   PM1<3> = PM1_3
*                   PM1<2> = PM1_2
*                   PM1<1> = PM1_1
*                   PM1<0> = PM1_0
*                   PM2<3> = PM2_3
*                   PM2<2> = PM2_2
*                   PM2<1> = PM2_1
*                   PM2<0> = PM2_0
*                   PM3<3> = PM3_3
*                   PM3<2> = PM3_2
*                   PM3<1> = PM3_1
*                   PM3<0> = PM3_0
*                   RESET = RESET
.SUBCKT PMSM_G32 CLK NPM0_3 NPM0_2 NPM0_1 NPM0_0 NPM1_3 NPM1_2 NPM1_1 NPM1_0 
+NPM2_3 NPM2_2 NPM2_1 NPM2_0 NPM3_3 NPM3_2 NPM3_1 NPM3_0 PM0_3 PM0_2 PM0_1 
+PM0_0 PM1_3 PM1_2 PM1_1 PM1_0 PM2_3 PM2_2 PM2_1 PM2_0 PM3_3 PM3_2 PM3_1 PM3_0 
+RESET 
XU193 N123 N124 N125 N17 N122 OAI22X1_G10 
XU248 N182 N183 N174 N180 NAND3X1_G11 
XU245 NPM3_3 NPM2_3 NPM1_3 N177 NAND3X1_G11 
XU218 N153 N154 N144 N151 NAND3X1_G11 
XU215 NPM2_3 NPM0_3 NPM3_3 N148 NAND3X1_G11 
XU196 NPM3_3 NPM0_3 N129 N128 NAND3X1_G11 
XU188 NPM3_3 N67 N2 N189_0_ NAND3X1_G11 
XU204 N135 N136 N17 N134 NAND3X1_G11 
XU205 N137 N89 NPM2_0 N135 NAND3X1_G11 
XU231 N166 NPM1_0 N167 N165 AOI21X1_G3 
XU192 N120 N121 N122 N119 AOI21X1_G3 
XU281 NPM3_1 N112 NPM3_0 N195 AOI21X1_G3 
XU270 N193 NPM0_0 N140 N192 AOI21X1_G3 
XU263 N191 NPM0_0 N171 N190 AOI21X1_G3 
XU240 N169 NPM1_0 N170 N168 AOI21X1_G3 
XU228 NPM3_1 N81 NPM3_0 N164 AOI21X1_G3 
XU202 NPM3_1 N28 NPM3_0 N133 AOI21X1_G3 
XNPM0NORM_REG_3_ N189_0_ NPM0NORM146_3_ NPM0NORM_3 LATCH_G12 
XNPM2NORM_REG_3_ N189_0_ NPM2NORM174_3_ NPM2NORM_3 LATCH_G12 
XNPM3NORM_REG_3_ N189_0_ NPM3NORM188_3_ NPM3NORM_3 LATCH_G12 
XNPM1NORM_REG_3_ N189_0_ NPM1NORM160_3_ NPM1NORM_3 LATCH_G12 
XNPM0NORM_REG_0_ N189_0_ NPM0NORM146_0_ NPM0NORM_0 LATCH_G12 
XNPM0NORM_REG_2_ N189_0_ NPM0NORM146_2_ NPM0NORM_2 LATCH_G12 
XNPM2NORM_REG_0_ N189_0_ NPM2NORM174_0_ NPM2NORM_0 LATCH_G12 
XNPM2NORM_REG_2_ N189_0_ NPM2NORM174_2_ NPM2NORM_2 LATCH_G12 
XNPM3NORM_REG_1_ N189_0_ NPM3NORM188_1_ NPM3NORM_1 LATCH_G12 
XNPM3NORM_REG_2_ N189_0_ NPM3NORM188_2_ NPM3NORM_2 LATCH_G12 
XNPM2NORM_REG_1_ N189_0_ NPM2NORM174_1_ NPM2NORM_1 LATCH_G12 
XNPM3NORM_REG_0_ N189_0_ NPM3NORM188_0_ NPM3NORM_0 LATCH_G12 
XNPM1NORM_REG_0_ N189_0_ NPM1NORM160_0_ NPM1NORM_0 LATCH_G12 
XNPM1NORM_REG_2_ N189_0_ NPM1NORM160_2_ NPM1NORM_2 LATCH_G12 
XNPM1NORM_REG_1_ N189_0_ NPM1NORM160_1_ NPM1NORM_1 LATCH_G12 
XNPM0NORM_REG_1_ N189_0_ NPM0NORM146_1_ NPM0NORM_1 LATCH_G12 
XU158 N95 N96 N94 XOR2X1_G2 
XU161 N99 NPM0_3 N95 XOR2X1_G2 
XU101 N38 N39 N37 XOR2X1_G2 
XU102 N40 NPM2_3 N39 XOR2X1_G2 
XU76 N4 N5 N3 XOR2X1_G2 
XU77 N6 NPM3_3 N5 XOR2X1_G2 
XU132 N64 N65 N63 XOR2X1_G2 
XU134 N68 NPM1_3 N64 XOR2X1_G2 
XU178 N112 N110 N114 XOR2X1_G2 
XU174 N114 N111 N113 XOR2X1_G2 
XU92 N24 N27 N26 XOR2X1_G2 
XU146 N84 N80 N83 XOR2X1_G2 
XU120 N52 NPM2_1 N57 XOR2X1_G2 
XU168 N101 NPM0_2 N106 XOR2X1_G2 
XU82 N16 N10 N15 XOR2X1_G2 
XU141 N70 NPM1_2 N75 XOR2X1_G2 
XU112 N17 N45 N50 XOR2X1_G2 
XU149 N81 N79 N84 XOR2X1_G2 
XU93 N21 NPM3_1 N27 XOR2X1_G2 
XU140 N73 N75 N74 XOR2X1_G2 
XU119 N55 N57 N56 XOR2X1_G2 
XU167 N104 N106 N105 XOR2X1_G2 
XU85 N19 N11 N16 XOR2X1_G2 
XU108 N50 N44 N49 XOR2X1_G2 
XU260 N181 N46 N184 N97 N189 AOI22X1_G1 
XU255 NPM0_2 N187 N188 N184 N186 AOI22X1_G1 
XU247 NPM0_2 N180 N181 N19 N179 AOI22X1_G1 
XU250 N184 N162 N185 N17 N178 AOI22X1_G1 
XU220 N155 N156 N157 N17 N149 AOI22X1_G1 
XU217 NPM1_2 N151 N152 N19 N150 AOI22X1_G1 
XU225 N152 N46 N155 N67 N161 AOI22X1_G1 
XU222 NPM1_2 N159 N120 N152 N158 AOI22X1_G1 
XU195 N127 N126 NPM2_3 N128 N118 AOI22X1_G1 
XU199 N19 N121 N121 NPM2_2 N131 AOI22X1_G1 
XU194 N121 N46 N126 N67 N125 AOI22X1_G1 
XU280 NPM0_1 N25 N195 NPM0_0 N194 AOI22X1_G1 
XU227 NPM1_1 N25 N164 NPM1_0 N163 AOI22X1_G1 
XU201 NPM2_1 N25 N133 NPM2_0 N132 AOI22X1_G1 
XU106 NPM0_3 N47 NPM1_3 N48 N14 AOI22X1_G1 
XU122 NPM0_1 N47 NPM1_1 N48 N29 AOI22X1_G1 
XU111 NPM0_2 N47 NPM1_2 N48 N18 AOI22X1_G1 
XU129 NPM0_0 N47 NPM1_0 N48 N35 AOI22X1_G1 
XU242 N172 N173 N47 NOR2X1_G7 
XU212 N142 N143 N48 NOR2X1_G7 
XU124 N59 N13 N36 NOR2X1_G7 
XU181 N87 N48 N93 NOR2X1_G7 
XU157 N93 N94 NPM0NORM146_3_ NOR2X1_G7 
XU100 N36 N37 NPM2NORM174_3_ NOR2X1_G7 
XU75 N2 N3 NPM3NORM188_3_ NOR2X1_G7 
XU265 NPM1_0 N170 N191 NOR2X1_G7 
XU241 NPM0_0 N171 N169 NOR2X1_G7 
XU271 N112 NPM2_1 N140 NOR2X1_G7 
XU264 N112 NPM1_1 N171 NOR2X1_G7 
XU266 N81 NPM0_1 N170 NOR2X1_G7 
XU211 N47 N48 N87 NOR2X1_G7 
XU152 N47 N87 N62 NOR2X1_G7 
XU131 N62 N63 NPM1NORM160_3_ NOR2X1_G7 
XU180 N115 N93 NPM0NORM146_0_ NOR2X1_G7 
XU173 N93 N113 NPM0NORM146_1_ NOR2X1_G7 
XU95 N30 N2 NPM3NORM188_0_ NOR2X1_G7 
XU151 N86 N62 NPM1NORM160_0_ NOR2X1_G7 
XU123 N58 N36 NPM2NORM174_0_ NOR2X1_G7 
XU189 N13 N98 N2 NOR2X1_G7 
XU81 N2 N15 NPM3NORM188_2_ NOR2X1_G7 
XU118 N36 N56 NPM2NORM174_1_ NOR2X1_G7 
XU107 N36 N49 NPM2NORM174_2_ NOR2X1_G7 
XU166 N93 N105 NPM0NORM146_2_ NOR2X1_G7 
XU139 N62 N74 NPM1NORM160_2_ NOR2X1_G7 
XU91 N2 N26 NPM3NORM188_1_ NOR2X1_G7 
XU145 N62 N83 NPM1NORM160_1_ NOR2X1_G7 
XU159 N97 N66 N48 N96 MUX2X1_G5 
XU133 N67 N66 N47 N65 MUX2X1_G5 
XU160 NPM2_3 NPM3_3 N98 N66 MUX2X1_G5 
XU171 NPM1_2 N82 N48 N104 MUX2X1_G5 
XU176 NPM1_1 N85 N48 N107 MUX2X1_G5 
XU177 N25 N28 N59 N85 MUX2X1_G5 
XU144 NPM0_2 N82 N47 N73 MUX2X1_G5 
XU148 NPM0_1 N85 N47 N76 MUX2X1_G5 
XU185 N89 N91 N48 N117 MUX2X1_G5 
XU186 NPM2_0 NPM3_0 N98 N91 MUX2X1_G5 
XU156 N92 N91 N47 N90 MUX2X1_G5 
XU172 N19 N17 N59 N82 MUX2X1_G5 
XU259 NPM2_3 N174 N189 N187 OAI21X1_G4 
XU254 N183 N160 N186 N172 OAI21X1_G4 
XU244 N176 N177 NPM0_3 N175 OAI21X1_G4 
XU243 N174 N145 N175 N173 OAI21X1_G4 
XU230 NPM2_2 N162 N165 N157 OAI21X1_G4 
XU224 NPM2_3 N144 N161 N159 OAI21X1_G4 
XU221 N153 N141 N158 N142 OAI21X1_G4 
XU213 N144 N145 N146 N143 OAI21X1_G4 
XU214 N147 N148 NPM1_3 N146 OAI21X1_G4 
XU198 N123 NPM1_2 N131 N130 OAI21X1_G4 
XU105 N46 N13 N14 N38 OAI21X1_G4 
XU80 N12 N13 N14 N4 OAI21X1_G4 
XU279 NPM3_2 N156 N194 N181 OAI21X1_G4 
XU269 NPM2_2 N156 N192 N185 OAI21X1_G4 
XU262 NPM1_2 N156 N190 N184 OAI21X1_G4 
XU239 NPM0_2 N162 N168 N155 OAI21X1_G4 
XU226 NPM3_2 N162 N163 N152 OAI21X1_G4 
XU200 NPM3_2 N17 N132 N121 OAI21X1_G4 
XU207 N34 N138 N139 N126 OAI21X1_G4 
XU136 N72 N73 NPM1_2 N71 OAI21X1_G4 
XU135 N69 N70 N71 N68 OAI21X1_G4 
XU183 N92 N117 N108 N116 OAI21X1_G4 
XU169 N107 N108 N109 N101 OAI21X1_G4 
XU170 N110 N111 N112 N109 OAI21X1_G4 
XU128 N13 N33 N35 N61 OAI21X1_G4 
XU154 N89 N90 N77 N88 OAI21X1_G4 
XU79 N10 N11 NPM3_2 N9 OAI21X1_G4 
XU103 N41 N42 N43 N40 OAI21X1_G4 
XU142 N76 N77 N78 N70 OAI21X1_G4 
XU114 N51 N52 N53 N42 OAI21X1_G4 
XU126 N34 N61 N52 N60 OAI21X1_G4 
XU163 N103 N104 NPM0_2 N102 OAI21X1_G4 
XU78 N7 N8 N9 N6 OAI21X1_G4 
XU121 N25 N13 N29 N55 OAI21X1_G4 
XU87 N20 N21 N22 N8 OAI21X1_G4 
XU104 N44 N45 NPM2_2 N43 OAI21X1_G4 
XU143 N79 N80 N81 N78 OAI21X1_G4 
XU99 N34 N13 N35 N32 OAI21X1_G4 
XU115 N54 N55 N28 N53 OAI21X1_G4 
XU162 N100 N101 N102 N99 OAI21X1_G4 
XU84 N17 N13 N18 N7 OAI21X1_G4 
XU94 N28 N13 N29 N24 OAI21X1_G4 
XU88 N23 N24 N25 N22 OAI21X1_G4 
XU110 N13 N19 N18 N41 OAI21X1_G4 
XU97 N32 N33 N21 N31 OAI21X1_G4 
XU246 N178 N179 N176 NAND2X1_G9 
XU216 N149 N150 N147 NAND2X1_G9 
XU191 N118 N119 N59 NAND2X1_G9 
XU275 N19 N46 N160 NAND2X1_G9 
XU273 NPM2_1 N112 N139 NAND2X1_G9 
XU257 N162 N97 N124 NAND2X1_G9 
XU251 N17 N12 N145 NAND2X1_G9 
XU237 N156 N67 N141 NAND2X1_G9 
XU236 NPM2_1 N81 N136 NAND2X1_G9 
XU233 NPM1_1 N28 N137 NAND2X1_G9 
XU98 N33 N32 N21 NAND2X1_G9 
XU127 N34 N61 N52 NAND2X1_G9 
XU155 N90 N89 N77 NAND2X1_G9 
XU184 N117 N92 N108 NAND2X1_G9 
XU256 N124 N188 INVX1_G6 
XU249 N184 N182 INVX1_G6 
XU232 N137 N167 INVX1_G6 
XU219 N152 N154 INVX1_G6 
XU209 N141 N127 INVX1_G6 
XU197 N130 N129 INVX1_G6 
XU203 N134 N123 INVX1_G6 
XU206 NPM1_0 N89 INVX1_G6 
XU276 NPM3_3 N46 INVX1_G6 
XU261 NPM1_3 N97 INVX1_G6 
XU285 NPM0_3 N67 INVX1_G6 
XU284 NPM0_2 N156 INVX1_G6 
XU283 NPM3_1 N25 INVX1_G6 
XU282 NPM0_1 N112 INVX1_G6 
XU278 N181 N183 INVX1_G6 
XU277 NPM3_2 N19 INVX1_G6 
XU223 N160 N120 INVX1_G6 
XU268 N185 N174 INVX1_G6 
XU274 NPM2_0 N34 INVX1_G6 
XU267 NPM1_1 N81 INVX1_G6 
XU258 NPM1_2 N162 INVX1_G6 
XU253 NPM2_2 N17 INVX1_G6 
XU252 NPM2_3 N12 INVX1_G6 
XU238 N155 N153 INVX1_G6 
XU229 N157 N144 INVX1_G6 
XU234 NPM2_1 N28 INVX1_G6 
XU210 N87 N13 INVX1_G6 
XU137 N70 N72 INVX1_G6 
XU138 N73 N69 INVX1_G6 
XU182 N116 N115 INVX1_G6 
XU175 N107 N111 INVX1_G6 
XU90 N24 N20 INVX1_G6 
XU153 N88 N86 INVX1_G6 
XU130 NPM3_0 N33 INVX1_G6 
XU150 N77 N79 INVX1_G6 
XU117 N55 N51 INVX1_G6 
XU165 N104 N100 INVX1_G6 
XU187 NPM0_0 N92 INVX1_G6 
XU83 N7 N10 INVX1_G6 
XU116 N52 N54 INVX1_G6 
XU125 N60 N58 INVX1_G6 
XU113 N42 N45 INVX1_G6 
XU89 N21 N23 INVX1_G6 
XU164 N101 N103 INVX1_G6 
XU179 N108 N110 INVX1_G6 
XU96 N31 N30 INVX1_G6 
XU109 N41 N44 INVX1_G6 
XU190 N59 N98 INVX1_G6 
XU74 RESET N1 INVX1_G6 
XU147 N76 N80 INVX1_G6 
XU86 N8 N11 INVX1_G6 
XU235 N34 N136 N166 AND2X1_G8 
XU272 N34 N139 N193 AND2X1_G8 
XU72 NPM0NORM_1 N1 PM0233_1_ AND2X1_G8 
XU71 NPM0NORM_2 N1 PM0233_2_ AND2X1_G8 
XU73 NPM0NORM_0 N1 PM0233_0_ AND2X1_G8 
XU70 NPM0NORM_3 N1 PM0233_3_ AND2X1_G8 
XU208 N140 NPM0_0 N138 OR2X1_G13 
XU61 NPM3NORM_0 RESET PM3254_0_ OR2X1_G13 
XU63 NPM2NORM_2 RESET PM2247_2_ OR2X1_G13 
XU65 NPM2NORM_0 RESET PM2247_0_ OR2X1_G13 
XU62 NPM2NORM_3 RESET PM2247_3_ OR2X1_G13 
XU64 NPM2NORM_1 RESET PM2247_1_ OR2X1_G13 
XU59 NPM3NORM_2 RESET PM3254_2_ OR2X1_G13 
XU67 NPM1NORM_2 RESET PM1240_2_ OR2X1_G13 
XU58 NPM3NORM_3 RESET PM3254_3_ OR2X1_G13 
XU69 NPM1NORM_0 RESET PM1240_0_ OR2X1_G13 
XU60 NPM3NORM_1 RESET PM3254_1_ OR2X1_G13 
XU66 NPM1NORM_3 RESET PM1240_3_ OR2X1_G13 
XU68 NPM1NORM_1 RESET PM1240_1_ OR2X1_G13 
XPM3_REG_3_ CLK PM3254_3_ PM3_3 DFFPOSX1_G14 
XPM3_REG_0_ CLK PM3254_0_ PM3_0 DFFPOSX1_G14 
XPM1_REG_2_ CLK PM1240_2_ PM1_2 DFFPOSX1_G14 
XPM2_REG_2_ CLK PM2247_2_ PM2_2 DFFPOSX1_G14 
XPM1_REG_3_ CLK PM1240_3_ PM1_3 DFFPOSX1_G14 
XPM0_REG_3_ CLK PM0233_3_ PM0_3 DFFPOSX1_G14 
XPM1_REG_1_ CLK PM1240_1_ PM1_1 DFFPOSX1_G14 
XPM3_REG_2_ CLK PM3254_2_ PM3_2 DFFPOSX1_G14 
XPM0_REG_0_ CLK PM0233_0_ PM0_0 DFFPOSX1_G14 
XPM0_REG_2_ CLK PM0233_2_ PM0_2 DFFPOSX1_G14 
XPM0_REG_1_ CLK PM0233_1_ PM0_1 DFFPOSX1_G14 
XPM1_REG_0_ CLK PM1240_0_ PM1_0 DFFPOSX1_G14 
XPM2_REG_0_ CLK PM2247_0_ PM2_0 DFFPOSX1_G14 
XPM2_REG_1_ CLK PM2247_1_ PM2_1 DFFPOSX1_G14 
XPM2_REG_3_ CLK PM2247_3_ PM2_3 DFFPOSX1_G14 
XPM3_REG_1_ CLK PM3254_1_ PM3_1 DFFPOSX1_G14 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS PMSM_G32 
* FILE NAME: OSU_STDCELLS_AOI22X1_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: AOI22X1.
* GENERATED FOR: HSPICES.
* GENERATED ON NOV  7 08:54:31 2007.
   
* TERMINAL MAPPING: A = A
*                   B = B
*                   C = C
*                   D = D
*                   Y = Y
.SUBCKT AOI22X1_G1 A B C D Y 
M23 Y B NET10 0  TSMC20N  L=200E-9 W=2E-6 AD=1E-12 AS=1E-12 PD=5E-6 PS=5E-6 
+M=1 
M24 NET10 A 0 0  TSMC20N  L=200E-9 W=2E-6 AD=1E-12 AS=1E-12 PD=5E-6 PS=5E-6 
+M=1 
M25 Y C NET037 0  TSMC20N  L=200E-9 W=2E-6 AD=1E-12 AS=1E-12 PD=5E-6 PS=5E-6 
+M=1 
M26 NET037 D 0 0  TSMC20N  L=200E-9 W=2E-6 AD=1E-12 AS=1E-12 PD=5E-6 PS=5E-6 
+M=1 
M19 NET22 A VDD! VDD!  TSMC20P  L=200E-9 W=4E-6 AD=2E-12 AS=2E-12 PD=9E-6 
+PS=9E-6 M=1 
M20 Y D NET22 VDD!  TSMC20P  L=200E-9 W=4E-6 AD=2E-12 AS=2E-12 PD=9E-6 PS=9E-6 
+M=1 
M21 NET22 B VDD! VDD!  TSMC20P  L=200E-9 W=4E-6 AD=2E-12 AS=2E-12 PD=9E-6 
+PS=9E-6 M=1 
M22 Y C NET22 VDD!  TSMC20P  L=200E-9 W=4E-6 AD=2E-12 AS=2E-12 PD=9E-6 PS=9E-6 
+M=1 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS AOI22X1_G1 
* FILE NAME: OSU_STDCELLS_XOR2X1_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: XOR2X1.
* GENERATED FOR: HSPICES.
* GENERATED ON NOV  7 08:54:31 2007.
   
* TERMINAL MAPPING: A = A
*                   B = B
*                   Y = Y
.SUBCKT XOR2X1_G2 A B Y 
M25 A_B A 0 0  TSMC20N  L=200E-9 W=2E-6 AD=1E-12 AS=1E-12 PD=5E-6 PS=5E-6 M=1 
M28 Y A_B NET12 0  TSMC20N  L=200E-9 W=2E-6 AD=1E-12 AS=1E-12 PD=5E-6 PS=5E-6 
+M=1 
M29 NET12 B_B 0 0  TSMC20N  L=200E-9 W=2E-6 AD=1E-12 AS=1E-12 PD=5E-6 PS=5E-6 
+M=1 
M30 NET9 B 0 0  TSMC20N  L=200E-9 W=2E-6 AD=1E-12 AS=1E-12 PD=5E-6 PS=5E-6 M=1 
M33 Y A NET9 0  TSMC20N  L=200E-9 W=2E-6 AD=1E-12 AS=1E-12 PD=5E-6 PS=5E-6 M=1 
M34 B_B B 0 0  TSMC20N  L=200E-9 W=2E-6 AD=1E-12 AS=1E-12 PD=5E-6 PS=5E-6 M=1 
M24 A_B A VDD! VDD!  TSMC20P  L=200E-9 W=4E-6 AD=2E-12 AS=2E-12 PD=9E-6 
+PS=9E-6 M=1 
M26 NET35 B_B VDD! VDD!  TSMC20P  L=200E-9 W=4E-6 AD=2E-12 AS=2E-12 PD=9E-6 
+PS=9E-6 M=1 
M27 Y A NET35 VDD!  TSMC20P  L=200E-9 W=4E-6 AD=2E-12 AS=2E-12 PD=9E-6 PS=9E-6 
+M=1 
M31 NET33 B VDD! VDD!  TSMC20P  L=200E-9 W=4E-6 AD=2E-12 AS=2E-12 PD=9E-6 
+PS=9E-6 M=1 
M32 Y A_B NET33 VDD!  TSMC20P  L=200E-9 W=4E-6 AD=2E-12 AS=2E-12 PD=9E-6 
+PS=9E-6 M=1 
M35 B_B B VDD! VDD!  TSMC20P  L=200E-9 W=4E-6 AD=2E-12 AS=2E-12 PD=9E-6 
+PS=9E-6 M=1 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS XOR2X1_G2 
* FILE NAME: OSU_STDCELLS_NAND2X1_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: NAND2X1.
* GENERATED FOR: HSPICES.
* GENERATED ON NOV  7 08:54:32 2007.
   
* TERMINAL MAPPING: A = A
*                   B = B
*                   Y = Y
.SUBCKT NAND2X1_G9 A B Y 
M9 Y A NET9 0  TSMC20N  L=200E-9 W=2E-6 AD=1E-12 AS=1E-12 PD=5E-6 PS=5E-6 M=1 
M12 NET9 B 0 0  TSMC20N  L=200E-9 W=2E-6 AD=1E-12 AS=1E-12 PD=5E-6 PS=5E-6 M=1 
M10 Y B VDD! VDD!  TSMC20P  L=200E-9 W=2E-6 AD=1E-12 AS=1E-12 PD=5E-6 PS=5E-6 
+M=1 
M11 Y A VDD! VDD!  TSMC20P  L=200E-9 W=2E-6 AD=1E-12 AS=1E-12 PD=5E-6 PS=5E-6 
+M=1 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS NAND2X1_G9 
* FILE NAME: VITERBI_SPDU_1_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: SPDU_1.
* GENERATED FOR: HSPICES.
* GENERATED ON NOV  7 08:54:34 2007.
   
* TERMINAL MAPPING: CLK = CLK
*                   D0 = D0
*                   D1 = D1
*                   D2 = D2
*                   D3 = D3
*                   IN0 = IN0
*                   IN1 = IN1
*                   IN2 = IN2
*                   IN3 = IN3
*                   OUT0 = OUT0
*                   OUT1 = OUT1
*                   OUT2 = OUT2
*                   OUT3 = OUT3
*                   RESET = RESET
.SUBCKT SPDU_1_G17 CLK D0 D1 D2 D3 IN0 IN1 IN2 IN3 OUT0 OUT1 OUT2 OUT3 RESET 
XOUT3_REG CLK OUT3223 OUT3 DFFPOSX1_G14 
XOUT2_REG CLK OUT2217 OUT2 DFFPOSX1_G14 
XOUT0_REG CLK OUT0205 OUT0 DFFPOSX1_G14 
XOUT1_REG CLK OUT1211 OUT1 DFFPOSX1_G14 
XU37 RESET N1 OUT3223 NOR2X1_G7 
XU43 RESET N4 OUT0205 NOR2X1_G7 
XU39 RESET N2 OUT2217 NOR2X1_G7 
XU41 RESET N3 OUT1211 NOR2X1_G7 
XU38 IN3 IN2 D3 N1 MUX2X1_G5 
XU44 IN1 IN0 D0 N4 MUX2X1_G5 
XU42 IN3 IN2 D1 N3 MUX2X1_G5 
XU40 IN1 IN0 D2 N2 MUX2X1_G5 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS SPDU_1_G17 
* FILE NAME: OSU_STDCELLS_MUX2X1_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: MUX2X1.
* GENERATED FOR: HSPICES.
* GENERATED ON NOV  7 08:54:31 2007.
   
* TERMINAL MAPPING: A = A
*                   B = B
*                   S = S
*                   Y = Y
.SUBCKT MUX2X1_G5 A B S Y 
M15 NET15 B VDD! VDD!  TSMC20P  L=200E-9 W=4E-6 AD=2E-12 AS=2E-12 PD=9E-6 
+PS=9E-6 M=1 
M16 S_B S VDD! VDD!  TSMC20P  L=200E-9 W=2E-6 AD=1E-12 AS=1E-12 PD=5E-6 
+PS=5E-6 M=1 
M17 Y S NET15 VDD!  TSMC20P  L=200E-9 W=4E-6 AD=2E-12 AS=2E-12 PD=9E-6 PS=9E-6 
+M=1 
M18 NET9 A VDD! VDD!  TSMC20P  L=200E-9 W=4E-6 AD=2E-12 AS=2E-12 PD=9E-6 
+PS=9E-6 M=1 
M19 Y S_B NET9 VDD!  TSMC20P  L=200E-9 W=4E-6 AD=2E-12 AS=2E-12 PD=9E-6 
+PS=9E-6 M=1 
M20 Y S_B NET34 0  TSMC20N  L=200E-9 W=2E-6 AD=1E-12 AS=1E-12 PD=5E-6 PS=5E-6 
+M=1 
M21 S_B S 0 0  TSMC20N  L=200E-9 W=1E-6 AD=500E-15 AS=500E-15 PD=3E-6 PS=3E-6 
+M=1 
M22 NET34 B 0 0  TSMC20N  L=200E-9 W=2E-6 AD=1E-12 AS=1E-12 PD=5E-6 PS=5E-6 
+M=1 
M23 Y S NET25 0  TSMC20N  L=200E-9 W=2E-6 AD=1E-12 AS=1E-12 PD=5E-6 PS=5E-6 
+M=1 
M24 NET25 A 0 0  TSMC20N  L=200E-9 W=2E-6 AD=1E-12 AS=1E-12 PD=5E-6 PS=5E-6 
+M=1 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS MUX2X1_G5 
* FILE NAME: OSU_STDCELLS_INVX1_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: INVX1.
* GENERATED FOR: HSPICES.
* GENERATED ON NOV  7 08:54:31 2007.
   
* TERMINAL MAPPING: A = A
*                   Y = Y
.SUBCKT INVX1_G6 A Y 
M4 Y A 0 0  TSMC20N  L=200E-9 W=1E-6 AD=500E-15 AS=500E-15 PD=3E-6 PS=3E-6 M=1 
M5 Y A VDD! VDD!  TSMC20P  L=200E-9 W=2E-6 AD=1E-12 AS=1E-12 PD=5E-6 PS=5E-6 
+M=1 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS INVX1_G6 
* FILE NAME: VITERBI_SELECTOR_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: SELECTOR.
* GENERATED FOR: HSPICES.
* GENERATED ON NOV  7 08:54:34 2007.
   
* TERMINAL MAPPING: D0 = D0
*                   D1 = D1
*                   PM0<3> = PM0_3
*                   PM0<2> = PM0_2
*                   PM0<1> = PM0_1
*                   PM0<0> = PM0_0
*                   PM1<3> = PM1_3
*                   PM1<2> = PM1_2
*                   PM1<1> = PM1_1
*                   PM1<0> = PM1_0
*                   PM2<3> = PM2_3
*                   PM2<2> = PM2_2
*                   PM2<1> = PM2_1
*                   PM2<0> = PM2_0
*                   PM3<3> = PM3_3
*                   PM3<2> = PM3_2
*                   PM3<1> = PM3_1
*                   PM3<0> = PM3_0
.SUBCKT SELECTOR_G16 D0 D1 PM0_3 PM0_2 PM0_1 PM0_0 PM1_3 PM1_2 PM1_1 PM1_0 
+PM2_3 PM2_2 PM2_1 PM2_0 PM3_3 PM3_2 PM3_1 PM3_0 
XU86 PM0_2 N16 PM0_1 N48 N44 OAI22X1_G10 
XU49 N13 N14 N15 N16 N12 OAI22X1_G10 
XU50 N13 N17 N15 N18 N11 OAI22X1_G10 
XU71 PM2_2 N31 PM2_1 N38 N33 OAI22X1_G10 
XU83 N46 PM0_2 PM0_3 N14 N45 AOI22X1_G1 
XU69 N35 PM2_2 PM2_3 N36 N34 AOI22X1_G1 
XU91 N50 N24 PM1_1 N49 OAI21X1_G4 
XU68 N32 N33 N34 N3 OAI21X1_G4 
XU82 N43 N44 N45 N2 OAI21X1_G4 
XU54 N19 N20 N21 N9 OAI21X1_G4 
XU77 N41 N42 PM3_1 N39 OAI21X1_G4 
XU47 N8 N9 N10 N7 OAI21X1_G4 
XU46 N5 N6 N7 N4 OAI21X1_G4 
XU56 N20 N19 N23 N22 AOI21X1_G3 
XU63 PM1_0 PM0_0 N2 N26 MUX2X1_G5 
XU64 N31 N30 N3 N8 MUX2X1_G5 
XU44 N3 N2 D1 N1 MUX2X1_G5 
XU61 N29 N28 N3 N27 MUX2X1_G5 
XU57 PM3_1 PM2_1 N3 N23 MUX2X1_G5 
XU66 N14 N17 N2 N6 MUX2X1_G5 
XU58 N25 N24 N2 N20 MUX2X1_G5 
XU48 N12 N11 N2 N10 MUX2X1_G5 
XU85 N16 N47 N46 AND2X1_G8 
XU52 N8 N9 N15 AND2X1_G8 
XU88 N49 N47 N43 NAND2X1_G9 
XU73 N39 N40 N32 NAND2X1_G9 
XU67 PM2_3 PM3_3 N5 NAND2X1_G9 
XU89 PM1_3 N17 N47 NAND2X1_G9 
XU80 N28 PM3_0 N38 NOR2X1_G7 
XU75 N36 PM2_3 N37 NOR2X1_G7 
XU70 PM3_2 N37 N35 NOR2X1_G7 
XU60 N26 N27 N19 NOR2X1_G7 
XU94 N51 PM1_0 N48 NOR2X1_G7 
XU93 N48 N50 INVX1_G6 
XU76 PM3_3 N36 INVX1_G6 
XU51 PM0_2 N18 INVX1_G6 
XU87 PM1_2 N16 INVX1_G6 
XU65 PM2_2 N30 INVX1_G6 
XU59 PM1_1 N25 INVX1_G6 
XU78 PM2_1 N42 INVX1_G6 
XU43 N1 D0 INVX1_G6 
XU74 N37 N40 INVX1_G6 
XU45 N4 D1 INVX1_G6 
XU55 N22 N21 INVX1_G6 
XU53 N5 N13 INVX1_G6 
XU90 PM0_3 N17 INVX1_G6 
XU84 PM1_3 N14 INVX1_G6 
XU95 PM0_0 N51 INVX1_G6 
XU62 PM3_0 N29 INVX1_G6 
XU92 PM0_1 N24 INVX1_G6 
XU81 PM2_0 N28 INVX1_G6 
XU72 PM3_2 N31 INVX1_G6 
XU79 N38 N41 INVX1_G6 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS SELECTOR_G16 
* FILE NAME: OSU_STDCELLS_NOR2X1_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: NOR2X1.
* GENERATED FOR: HSPICES.
* GENERATED ON NOV  7 08:54:32 2007.
   
* TERMINAL MAPPING: A = A
*                   B = B
*                   Y = Y
.SUBCKT NOR2X1_G7 A B Y 
M10 NET5 B VDD! VDD!  TSMC20P  L=200E-9 W=4E-6 AD=2E-12 AS=2E-12 PD=9E-6 
+PS=9E-6 M=1 
M11 Y A NET5 VDD!  TSMC20P  L=200E-9 W=4E-6 AD=2E-12 AS=2E-12 PD=9E-6 PS=9E-6 
+M=1 
M9 Y B 0 0  TSMC20N  L=200E-9 W=1E-6 AD=500E-15 AS=500E-15 PD=3E-6 PS=3E-6 M=1 
M12 Y A 0 0  TSMC20N  L=200E-9 W=1E-6 AD=500E-15 AS=500E-15 PD=3E-6 PS=3E-6 
+M=1 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS NOR2X1_G7 
* FILE NAME: VITERBI_SPDU_14_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: SPDU_14.
* GENERATED FOR: HSPICES.
* GENERATED ON NOV  7 08:54:35 2007.
   
* TERMINAL MAPPING: CLK = CLK
*                   D0 = D0
*                   D1 = D1
*                   D2 = D2
*                   D3 = D3
*                   IN0 = IN0
*                   IN1 = IN1
*                   IN2 = IN2
*                   IN3 = IN3
*                   OUT0 = OUT0
*                   OUT1 = OUT1
*                   OUT2 = OUT2
*                   OUT3 = OUT3
*                   RESET = RESET
.SUBCKT SPDU_14_G30 CLK D0 D1 D2 D3 IN0 IN1 IN2 IN3 OUT0 OUT1 OUT2 OUT3 RESET 
XOUT1_REG CLK OUT1211 OUT1 DFFPOSX1_G14 
XOUT0_REG CLK OUT0205 OUT0 DFFPOSX1_G14 
XOUT2_REG CLK OUT2217 OUT2 DFFPOSX1_G14 
XOUT3_REG CLK OUT3223 OUT3 DFFPOSX1_G14 
XU39 RESET N2 OUT2217 NOR2X1_G7 
XU41 RESET N3 OUT1211 NOR2X1_G7 
XU43 RESET N4 OUT0205 NOR2X1_G7 
XU37 RESET N1 OUT3223 NOR2X1_G7 
XU38 IN3 IN2 D3 N1 MUX2X1_G5 
XU40 IN1 IN0 D2 N2 MUX2X1_G5 
XU42 IN3 IN2 D1 N3 MUX2X1_G5 
XU44 IN1 IN0 D0 N4 MUX2X1_G5 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS SPDU_14_G30 
* FILE NAME: VITERBI_SPDU_7_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: SPDU_7.
* GENERATED FOR: HSPICES.
* GENERATED ON NOV  7 08:54:35 2007.
   
* TERMINAL MAPPING: CLK = CLK
*                   D0 = D0
*                   D1 = D1
*                   D2 = D2
*                   D3 = D3
*                   IN0 = IN0
*                   IN1 = IN1
*                   IN2 = IN2
*                   IN3 = IN3
*                   OUT0 = OUT0
*                   OUT1 = OUT1
*                   OUT2 = OUT2
*                   OUT3 = OUT3
*                   RESET = RESET
.SUBCKT SPDU_7_G23 CLK D0 D1 D2 D3 IN0 IN1 IN2 IN3 OUT0 OUT1 OUT2 OUT3 RESET 
XOUT0_REG CLK OUT0205 OUT0 DFFPOSX1_G14 
XOUT2_REG CLK OUT2217 OUT2 DFFPOSX1_G14 
XOUT1_REG CLK OUT1211 OUT1 DFFPOSX1_G14 
XOUT3_REG CLK OUT3223 OUT3 DFFPOSX1_G14 
XU37 RESET N1 OUT3223 NOR2X1_G7 
XU43 RESET N4 OUT0205 NOR2X1_G7 
XU39 RESET N2 OUT2217 NOR2X1_G7 
XU41 RESET N3 OUT1211 NOR2X1_G7 
XU38 IN3 IN2 D3 N1 MUX2X1_G5 
XU42 IN3 IN2 D1 N3 MUX2X1_G5 
XU44 IN1 IN0 D0 N4 MUX2X1_G5 
XU40 IN1 IN0 D2 N2 MUX2X1_G5 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS SPDU_7_G23 
* FILE NAME: VITERBI_ADD_COMPARE_SELECT_0_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: ADD_COMPARE_SELECT_0.
* GENERATED FOR: HSPICES.
* GENERATED ON NOV  7 08:54:32 2007.
   
* TERMINAL MAPPING: BM1<1> = BM1_1
*                   BM1<0> = BM1_0
*                   BM2<1> = BM2_1
*                   BM2<0> = BM2_0
*                   D = D
*                   NPM<3> = NPM_3
*                   NPM<2> = NPM_2
*                   NPM<1> = NPM_1
*                   NPM<0> = NPM_0
*                   PM1<3> = PM1_3
*                   PM1<2> = PM1_2
*                   PM1<1> = PM1_1
*                   PM1<0> = PM1_0
*                   PM2<3> = PM2_3
*                   PM2<2> = PM2_2
*                   PM2<1> = PM2_1
*                   PM2<0> = PM2_0
.SUBCKT SUB1 BM1_1 BM1_0 BM2_1 BM2_0 D NPM_3 NPM_2 NPM_1 NPM_0 PM1_3 PM1_2 
+PM1_1 PM1_0 PM2_3 PM2_2 PM2_1 PM2_0 
XU38 N17 N8 N6 N18 N16 AOI22X1_G1 
XU52 N32 N33 N31 XOR2X1_G2 
XU53 PM1_1 BM1_1 N33 XOR2X1_G2 
XU48 N29 N30 N28 XOR2X1_G2 
XU49 PM2_1 BM2_1 N30 XOR2X1_G2 
XU33 N9 N1 N10 D AOI21X1_G3 
XU43 N5 N19 N7 N17 AOI21X1_G3 
XU65 N26 BM1_1 PM1_1 N41 AOI21X1_G3 
XU64 N40 N32 N41 N36 AOI21X1_G3 
XU73 N22 BM2_1 PM2_1 N43 AOI21X1_G3 
XU72 N42 N29 N43 N39 AOI21X1_G3 
XU37 N3 N15 N16 N14 OAI21X1_G4 
XU36 N4 N13 N14 N12 OAI21X1_G4 
XU35 N1 N9 N12 N11 OAI21X1_G4 
XU45 N25 N26 N27 N24 OAI21X1_G4 
XU41 N21 N22 N23 N20 OAI21X1_G4 
XU59 N37 N38 N23 N15 OAI21X1_G4 
XU55 N34 N35 N27 N13 OAI21X1_G4 
XU32 N8 N7 D NPM_0 MUX2X1_G5 
XU31 N6 N5 D NPM_1 MUX2X1_G5 
XU30 N4 N3 D NPM_2 MUX2X1_G5 
XU29 N2 N1 D NPM_3 MUX2X1_G5 
XU34 N11 N10 INVX1_G6 
XU44 N24 N7 INVX1_G6 
XU50 N18 N5 INVX1_G6 
XU76 BM2_1 N42 INVX1_G6 
XU69 N2 N9 INVX1_G6 
XU40 N20 N8 INVX1_G6 
XU66 N32 N26 INVX1_G6 
XU54 N13 N3 INVX1_G6 
XU58 N15 N4 INVX1_G6 
XU39 N19 N6 INVX1_G6 
XU68 BM1_1 N40 INVX1_G6 
XU74 N29 N22 INVX1_G6 
XU46 PM1_0 BM1_0 N25 NOR2X1_G7 
XU42 PM2_0 BM2_0 N21 NOR2X1_G7 
XU57 PM1_2 N36 N34 NOR2X1_G7 
XU70 N38 PM2_3 N2 NOR2X1_G7 
XU62 N35 PM1_3 N1 NOR2X1_G7 
XU61 PM2_2 N39 N37 NOR2X1_G7 
XU63 PM1_2 N36 N35 AND2X1_G8 
XU71 PM2_2 N39 N38 AND2X1_G8 
XU51 N31 N27 N18 NAND2X1_G9 
XU47 N28 N23 N19 NAND2X1_G9 
XU56 PM1_3 N35 N27 NAND2X1_G9 
XU67 PM1_0 BM1_0 N32 NAND2X1_G9 
XU75 PM2_0 BM2_0 N29 NAND2X1_G9 
XU60 PM2_3 N38 N23 NAND2X1_G9 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS SUB1 
* FILE NAME: OSU_STDCELLS_OAI22X1_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: OAI22X1.
* GENERATED FOR: HSPICES.
* GENERATED ON NOV  7 08:54:33 2007.
   
* TERMINAL MAPPING: A = A
*                   B = B
*                   C = C
*                   D = D
*                   Y = Y
.SUBCKT OAI22X1_G10 A B C D Y 
M18 Y C NET029 0  TSMC20N  L=200E-9 W=2E-6 AD=1E-12 AS=1E-12 PD=5E-6 PS=5E-6 
+M=1 
M20 NET029 A 0 0  TSMC20N  L=200E-9 W=2E-6 AD=1E-12 AS=1E-12 PD=5E-6 PS=5E-6 
+M=1 
M21 NET029 B 0 0  TSMC20N  L=200E-9 W=2E-6 AD=1E-12 AS=1E-12 PD=5E-6 PS=5E-6 
+M=1 
M22 Y D NET029 0  TSMC20N  L=200E-9 W=2E-6 AD=1E-12 AS=1E-12 PD=5E-6 PS=5E-6 
+M=1 
M17 NET18 A VDD! VDD!  TSMC20P  L=200E-9 W=4E-6 AD=2E-12 AS=2E-12 PD=9E-6 
+PS=9E-6 M=1 
M19 Y B NET18 VDD!  TSMC20P  L=200E-9 W=4E-6 AD=2E-12 AS=2E-12 PD=9E-6 PS=9E-6 
+M=1 
M23 Y D NET053 VDD!  TSMC20P  L=200E-9 W=4E-6 AD=2E-12 AS=2E-12 PD=9E-6 
+PS=9E-6 M=1 
M24 NET053 C VDD! VDD!  TSMC20P  L=200E-9 W=4E-6 AD=2E-12 AS=2E-12 PD=9E-6 
+PS=9E-6 M=1 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS OAI22X1_G10 
* FILE NAME: OSU_STDCELLS_DFFPOSX1_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: DFFPOSX1.
* GENERATED FOR: HSPICES.
* GENERATED ON NOV  7 08:54:33 2007.
   
* TERMINAL MAPPING: CLK = CLK
*                   D = D
*                   Q = Q
.SUBCKT DFFPOSX1_G14 CLK D Q 
M64 NET071 NET33 0 0  TSMC20N  L=200E-9 W=1E-6 AD=500E-15 AS=500E-15 PD=3E-6 
+PS=3E-6 M=1 
M58 NET33 CLK NET18 0  TSMC20N  L=200E-9 W=1E-6 AD=500E-15 AS=500E-15 PD=3E-6 
+PS=3E-6 M=1 
M57 CLK_B CLK 0 0  TSMC20N  L=200E-9 W=2E-6 AD=1E-12 AS=1E-12 PD=5E-6 PS=5E-6 
+M=1 
M61 NET18 NET071 0 0  TSMC20N  L=200E-9 W=1E-6 AD=500E-15 AS=500E-15 PD=3E-6 
+PS=3E-6 M=1 
M60 Q NET27 0 0  TSMC20N  L=200E-9 W=2E-6 AD=1E-12 AS=1E-12 PD=5E-6 PS=5E-6 
+M=1 
M66 NET24 NET071 0 0  TSMC20N  L=200E-9 W=1E-6 AD=500E-15 AS=500E-15 PD=3E-6 
+PS=3E-6 M=1 
M65 NET27 CLK NET24 0  TSMC20N  L=200E-9 W=1E-6 AD=500E-15 AS=500E-15 PD=3E-6 
+PS=3E-6 M=1 
M67 NET9 Q 0 0  TSMC20N  L=200E-9 W=1E-6 AD=500E-15 AS=500E-15 PD=3E-6 PS=3E-6 
+M=1 
M62 NET33 CLK_B NET30 0  TSMC20N  L=200E-9 W=1E-6 AD=500E-15 AS=500E-15 
+PD=3E-6 PS=3E-6 M=1 
M59 NET27 CLK_B NET9 0  TSMC20N  L=200E-9 W=1E-6 AD=500E-15 AS=500E-15 PD=3E-6 
+PS=3E-6 M=1 
M63 NET30 D 0 0  TSMC20N  L=200E-9 W=1E-6 AD=500E-15 AS=500E-15 PD=3E-6 
+PS=3E-6 M=1 
M46 CLK_B CLK VDD! VDD!  TSMC20P  L=200E-9 W=4E-6 AD=2E-12 AS=2E-12 PD=9E-6 
+PS=9E-6 M=1 
M47 NET50 NET071 VDD! VDD!  TSMC20P  L=200E-9 W=2E-6 AD=1E-12 AS=1E-12 PD=5E-6 
+PS=5E-6 M=1 
M48 NET41 Q VDD! VDD!  TSMC20P  L=200E-9 W=1E-6 AD=500E-15 AS=500E-15 PD=3E-6 
+PS=3E-6 M=1 
M49 Q NET27 VDD! VDD!  TSMC20P  L=200E-9 W=4E-6 AD=2E-12 AS=2E-12 PD=9E-6 
+PS=9E-6 M=1 
M50 NET33 CLK_B NET50 VDD!  TSMC20P  L=200E-9 W=2E-6 AD=1E-12 AS=1E-12 PD=5E-6 
+PS=5E-6 M=1 
M51 NET62 D VDD! VDD!  TSMC20P  L=200E-9 W=2E-6 AD=1E-12 AS=1E-12 PD=5E-6 
+PS=5E-6 M=1 
M52 NET33 CLK NET62 VDD!  TSMC20P  L=200E-9 W=2E-6 AD=1E-12 AS=1E-12 PD=5E-6 
+PS=5E-6 M=1 
M53 NET56 NET071 VDD! VDD!  TSMC20P  L=200E-9 W=2E-6 AD=1E-12 AS=1E-12 PD=5E-6 
+PS=5E-6 M=1 
M54 NET27 CLK_B NET56 VDD!  TSMC20P  L=200E-9 W=2E-6 AD=1E-12 AS=1E-12 PD=5E-6 
+PS=5E-6 M=1 
M55 NET071 NET33 VDD! VDD!  TSMC20P  L=200E-9 W=2E-6 AD=1E-12 AS=1E-12 PD=5E-6 
+PS=5E-6 M=1 
M56 NET27 CLK NET41 VDD!  TSMC20P  L=200E-9 W=1E-6 AD=500E-15 AS=500E-15 
+PD=3E-6 PS=3E-6 M=1 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS DFFPOSX1_G14 
* FILE NAME: VITERBI_ADD_COMPARE_SELECT_1_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: ADD_COMPARE_SELECT_1.
* GENERATED FOR: HSPICES.
* GENERATED ON NOV  7 08:54:32 2007.
   
* TERMINAL MAPPING: BM1<1> = BM1_1
*                   BM1<0> = BM1_0
*                   BM2<1> = BM2_1
*                   BM2<0> = BM2_0
*                   D = D
*                   NPM<3> = NPM_3
*                   NPM<2> = NPM_2
*                   NPM<1> = NPM_1
*                   NPM<0> = NPM_0
*                   PM1<3> = PM1_3
*                   PM1<2> = PM1_2
*                   PM1<1> = PM1_1
*                   PM1<0> = PM1_0
*                   PM2<3> = PM2_3
*                   PM2<2> = PM2_2
*                   PM2<1> = PM2_1
*                   PM2<0> = PM2_0
.SUBCKT SUB3 BM1_1 BM1_0 BM2_1 BM2_0 D NPM_3 NPM_2 NPM_1 NPM_0 PM1_3 PM1_2 
+PM1_1 PM1_0 PM2_3 PM2_2 PM2_1 PM2_0 
XU38 N17 N8 N6 N18 N16 AOI22X1_G1 
XU52 N32 N33 N31 XOR2X1_G2 
XU53 PM1_1 BM1_1 N33 XOR2X1_G2 
XU48 N29 N30 N28 XOR2X1_G2 
XU49 PM2_1 BM2_1 N30 XOR2X1_G2 
XU33 N9 N1 N10 D AOI21X1_G3 
XU43 N5 N19 N7 N17 AOI21X1_G3 
XU65 N26 BM1_1 PM1_1 N41 AOI21X1_G3 
XU64 N40 N32 N41 N36 AOI21X1_G3 
XU72 N42 N29 N43 N39 AOI21X1_G3 
XU73 N22 BM2_1 PM2_1 N43 AOI21X1_G3 
XU37 N3 N15 N16 N14 OAI21X1_G4 
XU36 N4 N13 N14 N12 OAI21X1_G4 
XU35 N1 N9 N12 N11 OAI21X1_G4 
XU45 N25 N26 N27 N24 OAI21X1_G4 
XU41 N21 N22 N23 N20 OAI21X1_G4 
XU55 N34 N35 N27 N13 OAI21X1_G4 
XU59 N37 N38 N23 N15 OAI21X1_G4 
XU31 N6 N5 D NPM_1 MUX2X1_G5 
XU30 N4 N3 D NPM_2 MUX2X1_G5 
XU29 N2 N1 D NPM_3 MUX2X1_G5 
XU32 N8 N7 D NPM_0 MUX2X1_G5 
XU34 N11 N10 INVX1_G6 
XU44 N24 N7 INVX1_G6 
XU40 N20 N8 INVX1_G6 
XU76 BM2_1 N42 INVX1_G6 
XU54 N13 N3 INVX1_G6 
XU74 N29 N22 INVX1_G6 
XU68 BM1_1 N40 INVX1_G6 
XU39 N19 N6 INVX1_G6 
XU66 N32 N26 INVX1_G6 
XU50 N18 N5 INVX1_G6 
XU58 N15 N4 INVX1_G6 
XU69 N2 N9 INVX1_G6 
XU46 PM1_0 BM1_0 N25 NOR2X1_G7 
XU42 PM2_0 BM2_0 N21 NOR2X1_G7 
XU62 N35 PM1_3 N1 NOR2X1_G7 
XU70 N38 PM2_3 N2 NOR2X1_G7 
XU61 PM2_2 N39 N37 NOR2X1_G7 
XU57 PM1_2 N36 N34 NOR2X1_G7 
XU63 PM1_2 N36 N35 AND2X1_G8 
XU71 PM2_2 N39 N38 AND2X1_G8 
XU51 N31 N27 N18 NAND2X1_G9 
XU47 N28 N23 N19 NAND2X1_G9 
XU56 PM1_3 N35 N27 NAND2X1_G9 
XU60 PM2_3 N38 N23 NAND2X1_G9 
XU75 PM2_0 BM2_0 N29 NAND2X1_G9 
XU67 PM1_0 BM1_0 N32 NAND2X1_G9 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS SUB3 
* FILE NAME: OSU_STDCELLS_OAI21X1_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: OAI21X1.
* GENERATED FOR: HSPICES.
* GENERATED ON NOV  7 08:54:31 2007.
   
* TERMINAL MAPPING: A = A
*                   B = B
*                   C = C
*                   Y = Y
.SUBCKT OAI21X1_G4 A B C Y 
M15 Y C NET10 0  TSMC20N  L=200E-9 W=2E-6 AD=1E-12 AS=1E-12 PD=5E-6 PS=5E-6 
+M=1 
M19 NET10 A 0 0  TSMC20N  L=200E-9 W=2E-6 AD=1E-12 AS=1E-12 PD=5E-6 PS=5E-6 
+M=1 
M20 NET10 B 0 0  TSMC20N  L=200E-9 W=2E-6 AD=1E-12 AS=1E-12 PD=5E-6 PS=5E-6 
+M=1 
M16 NET18 A VDD! VDD!  TSMC20P  L=200E-9 W=4E-6 AD=2E-12 AS=2E-12 PD=9E-6 
+PS=9E-6 M=1 
M17 Y C VDD! VDD!  TSMC20P  L=200E-9 W=2E-6 AD=1E-12 AS=1E-12 PD=5E-6 PS=5E-6 
+M=1 
M18 Y B NET18 VDD!  TSMC20P  L=200E-9 W=4E-6 AD=2E-12 AS=2E-12 PD=9E-6 PS=9E-6 
+M=1 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS OAI21X1_G4 
* FILE NAME: VITERBI_ADD_COMPARE_SELECT_2_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: ADD_COMPARE_SELECT_2.
* GENERATED FOR: HSPICES.
* GENERATED ON NOV  7 08:54:32 2007.
   
* TERMINAL MAPPING: BM1<1> = BM1_1
*                   BM1<0> = BM1_0
*                   BM2<1> = BM2_1
*                   BM2<0> = BM2_0
*                   D = D
*                   NPM<3> = NPM_3
*                   NPM<2> = NPM_2
*                   NPM<1> = NPM_1
*                   NPM<0> = NPM_0
*                   PM1<3> = PM1_3
*                   PM1<2> = PM1_2
*                   PM1<1> = PM1_1
*                   PM1<0> = PM1_0
*                   PM2<3> = PM2_3
*                   PM2<2> = PM2_2
*                   PM2<1> = PM2_1
*                   PM2<0> = PM2_0
.SUBCKT SUB2 BM1_1 BM1_0 BM2_1 BM2_0 D NPM_3 NPM_2 NPM_1 NPM_0 PM1_3 PM1_2 
+PM1_1 PM1_0 PM2_3 PM2_2 PM2_1 PM2_0 
XU38 N17 N8 N6 N18 N16 AOI22X1_G1 
XU52 N32 N33 N31 XOR2X1_G2 
XU53 PM1_1 BM1_1 N33 XOR2X1_G2 
XU48 N29 N30 N28 XOR2X1_G2 
XU49 PM2_1 BM2_1 N30 XOR2X1_G2 
XU33 N9 N1 N10 D AOI21X1_G3 
XU43 N5 N19 N7 N17 AOI21X1_G3 
XU73 N22 BM2_1 PM2_1 N43 AOI21X1_G3 
XU72 N42 N29 N43 N39 AOI21X1_G3 
XU65 N26 BM1_1 PM1_1 N41 AOI21X1_G3 
XU64 N40 N32 N41 N36 AOI21X1_G3 
XU37 N3 N15 N16 N14 OAI21X1_G4 
XU36 N4 N13 N14 N12 OAI21X1_G4 
XU35 N1 N9 N12 N11 OAI21X1_G4 
XU45 N25 N26 N27 N24 OAI21X1_G4 
XU55 N34 N35 N27 N13 OAI21X1_G4 
XU59 N37 N38 N23 N15 OAI21X1_G4 
XU41 N21 N22 N23 N20 OAI21X1_G4 
XU31 N6 N5 D NPM_1 MUX2X1_G5 
XU30 N4 N3 D NPM_2 MUX2X1_G5 
XU29 N2 N1 D NPM_3 MUX2X1_G5 
XU32 N8 N7 D NPM_0 MUX2X1_G5 
XU34 N11 N10 INVX1_G6 
XU44 N24 N7 INVX1_G6 
XU66 N32 N26 INVX1_G6 
XU58 N15 N4 INVX1_G6 
XU54 N13 N3 INVX1_G6 
XU74 N29 N22 INVX1_G6 
XU39 N19 N6 INVX1_G6 
XU68 BM1_1 N40 INVX1_G6 
XU69 N2 N9 INVX1_G6 
XU50 N18 N5 INVX1_G6 
XU40 N20 N8 INVX1_G6 
XU76 BM2_1 N42 INVX1_G6 
XU46 PM1_0 BM1_0 N25 NOR2X1_G7 
XU62 N35 PM1_3 N1 NOR2X1_G7 
XU61 PM2_2 N39 N37 NOR2X1_G7 
XU42 PM2_0 BM2_0 N21 NOR2X1_G7 
XU57 PM1_2 N36 N34 NOR2X1_G7 
XU70 N38 PM2_3 N2 NOR2X1_G7 
XU71 PM2_2 N39 N38 AND2X1_G8 
XU63 PM1_2 N36 N35 AND2X1_G8 
XU51 N31 N27 N18 NAND2X1_G9 
XU47 N28 N23 N19 NAND2X1_G9 
XU56 PM1_3 N35 N27 NAND2X1_G9 
XU60 PM2_3 N38 N23 NAND2X1_G9 
XU75 PM2_0 BM2_0 N29 NAND2X1_G9 
XU67 PM1_0 BM1_0 N32 NAND2X1_G9 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS SUB2 
* FILE NAME: VITERBI_SPDU_8_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: SPDU_8.
* GENERATED FOR: HSPICES.
* GENERATED ON NOV  7 08:54:35 2007.
   
* TERMINAL MAPPING: CLK = CLK
*                   D0 = D0
*                   D1 = D1
*                   D2 = D2
*                   D3 = D3
*                   IN0 = IN0
*                   IN1 = IN1
*                   IN2 = IN2
*                   IN3 = IN3
*                   OUT0 = OUT0
*                   OUT1 = OUT1
*                   OUT2 = OUT2
*                   OUT3 = OUT3
*                   RESET = RESET
.SUBCKT SPDU_8_G24 CLK D0 D1 D2 D3 IN0 IN1 IN2 IN3 OUT0 OUT1 OUT2 OUT3 RESET 
XOUT2_REG CLK OUT2217 OUT2 DFFPOSX1_G14 
XOUT3_REG CLK OUT3223 OUT3 DFFPOSX1_G14 
XOUT1_REG CLK OUT1211 OUT1 DFFPOSX1_G14 
XOUT0_REG CLK OUT0205 OUT0 DFFPOSX1_G14 
XU37 RESET N1 OUT3223 NOR2X1_G7 
XU43 RESET N4 OUT0205 NOR2X1_G7 
XU39 RESET N2 OUT2217 NOR2X1_G7 
XU41 RESET N3 OUT1211 NOR2X1_G7 
XU38 IN3 IN2 D3 N1 MUX2X1_G5 
XU40 IN1 IN0 D2 N2 MUX2X1_G5 
XU44 IN1 IN0 D0 N4 MUX2X1_G5 
XU42 IN3 IN2 D1 N3 MUX2X1_G5 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS SPDU_8_G24 
* FILE NAME: VITERBI_SPDU_13_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: SPDU_13.
* GENERATED FOR: HSPICES.
* GENERATED ON NOV  7 08:54:35 2007.
   
* TERMINAL MAPPING: CLK = CLK
*                   D0 = D0
*                   D1 = D1
*                   D2 = D2
*                   D3 = D3
*                   IN0 = IN0
*                   IN1 = IN1
*                   IN2 = IN2
*                   IN3 = IN3
*                   OUT0 = OUT0
*                   OUT1 = OUT1
*                   OUT2 = OUT2
*                   OUT3 = OUT3
*                   RESET = RESET
.SUBCKT SPDU_13_G29 CLK D0 D1 D2 D3 IN0 IN1 IN2 IN3 OUT0 OUT1 OUT2 OUT3 RESET 
XOUT2_REG CLK OUT2217 OUT2 DFFPOSX1_G14 
XOUT3_REG CLK OUT3223 OUT3 DFFPOSX1_G14 
XOUT0_REG CLK OUT0205 OUT0 DFFPOSX1_G14 
XOUT1_REG CLK OUT1211 OUT1 DFFPOSX1_G14 
XU43 RESET N4 OUT0205 NOR2X1_G7 
XU37 RESET N1 OUT3223 NOR2X1_G7 
XU41 RESET N3 OUT1211 NOR2X1_G7 
XU39 RESET N2 OUT2217 NOR2X1_G7 
XU38 IN3 IN2 D3 N1 MUX2X1_G5 
XU44 IN1 IN0 D0 N4 MUX2X1_G5 
XU42 IN3 IN2 D1 N3 MUX2X1_G5 
XU40 IN1 IN0 D2 N2 MUX2X1_G5 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS SPDU_13_G29 
* FILE NAME: VITERBI_SPDU_11_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: SPDU_11.
* GENERATED FOR: HSPICES.
* GENERATED ON NOV  7 08:54:35 2007.
   
* TERMINAL MAPPING: CLK = CLK
*                   D0 = D0
*                   D1 = D1
*                   D2 = D2
*                   D3 = D3
*                   IN0 = IN0
*                   IN1 = IN1
*                   IN2 = IN2
*                   IN3 = IN3
*                   OUT0 = OUT0
*                   OUT1 = OUT1
*                   OUT2 = OUT2
*                   OUT3 = OUT3
*                   RESET = RESET
.SUBCKT SPDU_11_G27 CLK D0 D1 D2 D3 IN0 IN1 IN2 IN3 OUT0 OUT1 OUT2 OUT3 RESET 
XOUT3_REG CLK OUT3223 OUT3 DFFPOSX1_G14 
XOUT0_REG CLK OUT0205 OUT0 DFFPOSX1_G14 
XOUT1_REG CLK OUT1211 OUT1 DFFPOSX1_G14 
XOUT2_REG CLK OUT2217 OUT2 DFFPOSX1_G14 
XU39 RESET N2 OUT2217 NOR2X1_G7 
XU37 RESET N1 OUT3223 NOR2X1_G7 
XU43 RESET N4 OUT0205 NOR2X1_G7 
XU41 RESET N3 OUT1211 NOR2X1_G7 
XU38 IN3 IN2 D3 N1 MUX2X1_G5 
XU44 IN1 IN0 D0 N4 MUX2X1_G5 
XU40 IN1 IN0 D2 N2 MUX2X1_G5 
XU42 IN3 IN2 D1 N3 MUX2X1_G5 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS SPDU_11_G27 
* FILE NAME: VITERBI_SPDU_4_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: SPDU_4.
* GENERATED FOR: HSPICES.
* GENERATED ON NOV  7 08:54:34 2007.
   
* TERMINAL MAPPING: CLK = CLK
*                   D0 = D0
*                   D1 = D1
*                   D2 = D2
*                   D3 = D3
*                   IN0 = IN0
*                   IN1 = IN1
*                   IN2 = IN2
*                   IN3 = IN3
*                   OUT0 = OUT0
*                   OUT1 = OUT1
*                   OUT2 = OUT2
*                   OUT3 = OUT3
*                   RESET = RESET
.SUBCKT SPDU_4_G20 CLK D0 D1 D2 D3 IN0 IN1 IN2 IN3 OUT0 OUT1 OUT2 OUT3 RESET 
XOUT2_REG CLK OUT2217 OUT2 DFFPOSX1_G14 
XOUT1_REG CLK OUT1211 OUT1 DFFPOSX1_G14 
XOUT3_REG CLK OUT3223 OUT3 DFFPOSX1_G14 
XOUT0_REG CLK OUT0205 OUT0 DFFPOSX1_G14 
XU43 RESET N4 OUT0205 NOR2X1_G7 
XU37 RESET N1 OUT3223 NOR2X1_G7 
XU41 RESET N3 OUT1211 NOR2X1_G7 
XU39 RESET N2 OUT2217 NOR2X1_G7 
XU38 IN3 IN2 D3 N1 MUX2X1_G5 
XU40 IN1 IN0 D2 N2 MUX2X1_G5 
XU44 IN1 IN0 D0 N4 MUX2X1_G5 
XU42 IN3 IN2 D1 N3 MUX2X1_G5 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS SPDU_4_G20 
* FILE NAME: VITERBI_ADD_COMPARE_SELECT_3_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: ADD_COMPARE_SELECT_3.
* GENERATED FOR: HSPICES.
* GENERATED ON NOV  7 08:54:32 2007.
   
* TERMINAL MAPPING: BM1<1> = BM1_1
*                   BM1<0> = BM1_0
*                   BM2<1> = BM2_1
*                   BM2<0> = BM2_0
*                   D = D
*                   NPM<3> = NPM_3
*                   NPM<2> = NPM_2
*                   NPM<1> = NPM_1
*                   NPM<0> = NPM_0
*                   PM1<3> = PM1_3
*                   PM1<2> = PM1_2
*                   PM1<1> = PM1_1
*                   PM1<0> = PM1_0
*                   PM2<3> = PM2_3
*                   PM2<2> = PM2_2
*                   PM2<1> = PM2_1
*                   PM2<0> = PM2_0
.SUBCKT SUB4 BM1_1 BM1_0 BM2_1 BM2_0 D NPM_3 NPM_2 NPM_1 NPM_0 PM1_3 PM1_2 
+PM1_1 PM1_0 PM2_3 PM2_2 PM2_1 PM2_0 
XU38 N17 N8 N6 N18 N16 AOI22X1_G1 
XU52 N32 N33 N31 XOR2X1_G2 
XU53 PM1_1 BM1_1 N33 XOR2X1_G2 
XU48 N29 N30 N28 XOR2X1_G2 
XU49 PM2_1 BM2_1 N30 XOR2X1_G2 
XU33 N9 N1 N10 D AOI21X1_G3 
XU43 N5 N19 N7 N17 AOI21X1_G3 
XU73 N22 BM2_1 PM2_1 N43 AOI21X1_G3 
XU72 N42 N29 N43 N39 AOI21X1_G3 
XU65 N26 BM1_1 PM1_1 N41 AOI21X1_G3 
XU64 N40 N32 N41 N36 AOI21X1_G3 
XU37 N3 N15 N16 N14 OAI21X1_G4 
XU36 N4 N13 N14 N12 OAI21X1_G4 
XU35 N1 N9 N12 N11 OAI21X1_G4 
XU45 N25 N26 N27 N24 OAI21X1_G4 
XU55 N34 N35 N27 N13 OAI21X1_G4 
XU59 N37 N38 N23 N15 OAI21X1_G4 
XU41 N21 N22 N23 N20 OAI21X1_G4 
XU30 N4 N3 D NPM_2 MUX2X1_G5 
XU31 N6 N5 D NPM_1 MUX2X1_G5 
XU32 N8 N7 D NPM_0 MUX2X1_G5 
XU29 N2 N1 D NPM_3 MUX2X1_G5 
XU34 N11 N10 INVX1_G6 
XU44 N24 N7 INVX1_G6 
XU40 N20 N8 INVX1_G6 
XU69 N2 N9 INVX1_G6 
XU50 N18 N5 INVX1_G6 
XU68 BM1_1 N40 INVX1_G6 
XU39 N19 N6 INVX1_G6 
XU58 N15 N4 INVX1_G6 
XU54 N13 N3 INVX1_G6 
XU66 N32 N26 INVX1_G6 
XU74 N29 N22 INVX1_G6 
XU76 BM2_1 N42 INVX1_G6 
XU46 PM1_0 BM1_0 N25 NOR2X1_G7 
XU62 N35 PM1_3 N1 NOR2X1_G7 
XU61 PM2_2 N39 N37 NOR2X1_G7 
XU70 N38 PM2_3 N2 NOR2X1_G7 
XU42 PM2_0 BM2_0 N21 NOR2X1_G7 
XU57 PM1_2 N36 N34 NOR2X1_G7 
XU63 PM1_2 N36 N35 AND2X1_G8 
XU71 PM2_2 N39 N38 AND2X1_G8 
XU51 N31 N27 N18 NAND2X1_G9 
XU47 N28 N23 N19 NAND2X1_G9 
XU56 PM1_3 N35 N27 NAND2X1_G9 
XU60 PM2_3 N38 N23 NAND2X1_G9 
XU75 PM2_0 BM2_0 N29 NAND2X1_G9 
XU67 PM1_0 BM1_0 N32 NAND2X1_G9 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS SUB4 
* FILE NAME: VITERBI_SPDU_9_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: SPDU_9.
* GENERATED FOR: HSPICES.
* GENERATED ON NOV  7 08:54:35 2007.
   
* TERMINAL MAPPING: CLK = CLK
*                   D0 = D0
*                   D1 = D1
*                   D2 = D2
*                   D3 = D3
*                   IN0 = IN0
*                   IN1 = IN1
*                   IN2 = IN2
*                   IN3 = IN3
*                   OUT0 = OUT0
*                   OUT1 = OUT1
*                   OUT2 = OUT2
*                   OUT3 = OUT3
*                   RESET = RESET
.SUBCKT SPDU_9_G25 CLK D0 D1 D2 D3 IN0 IN1 IN2 IN3 OUT0 OUT1 OUT2 OUT3 RESET 
XOUT1_REG CLK OUT1211 OUT1 DFFPOSX1_G14 
XOUT3_REG CLK OUT3223 OUT3 DFFPOSX1_G14 
XOUT2_REG CLK OUT2217 OUT2 DFFPOSX1_G14 
XOUT0_REG CLK OUT0205 OUT0 DFFPOSX1_G14 
XU39 RESET N2 OUT2217 NOR2X1_G7 
XU41 RESET N3 OUT1211 NOR2X1_G7 
XU37 RESET N1 OUT3223 NOR2X1_G7 
XU43 RESET N4 OUT0205 NOR2X1_G7 
XU38 IN3 IN2 D3 N1 MUX2X1_G5 
XU44 IN1 IN0 D0 N4 MUX2X1_G5 
XU40 IN1 IN0 D2 N2 MUX2X1_G5 
XU42 IN3 IN2 D1 N3 MUX2X1_G5 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS SPDU_9_G25 
* FILE NAME: VITERBI_SPDU_0_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: SPDU_0.
* GENERATED FOR: HSPICES.
* GENERATED ON NOV  7 08:54:34 2007.
   
* TERMINAL MAPPING: CLK = CLK
*                   D0 = D0
*                   D1 = D1
*                   D2 = D2
*                   D3 = D3
*                   IN0 = IN0
*                   IN1 = IN1
*                   IN2 = IN2
*                   IN3 = IN3
*                   OUT0 = OUT0
*                   OUT1 = OUT1
*                   OUT2 = OUT2
*                   OUT3 = OUT3
*                   RESET = RESET
.SUBCKT SPDU_0_G21 CLK D0 D1 D2 D3 IN0 IN1 IN2 IN3 OUT0 OUT1 OUT2 OUT3 RESET 
XOUT2_REG CLK OUT2217 OUT2 DFFPOSX1_G14 
XOUT1_REG CLK OUT1211 OUT1 DFFPOSX1_G14 
XOUT0_REG CLK OUT0205 OUT0 DFFPOSX1_G14 
XOUT3_REG CLK OUT3223 OUT3 DFFPOSX1_G14 
XU39 RESET N2 OUT2217 NOR2X1_G7 
XU43 RESET N4 OUT0205 NOR2X1_G7 
XU41 RESET N3 OUT1211 NOR2X1_G7 
XU37 RESET N1 OUT3223 NOR2X1_G7 
XU38 IN3 IN2 D3 N1 MUX2X1_G5 
XU40 IN1 IN0 D2 N2 MUX2X1_G5 
XU42 IN3 IN2 D1 N3 MUX2X1_G5 
XU44 IN1 IN0 D0 N4 MUX2X1_G5 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS SPDU_0_G21 
* FILE NAME: OSU_STDCELLS_AOI21X1_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: AOI21X1.
* GENERATED FOR: HSPICES.
* GENERATED ON NOV  7 08:54:31 2007.
   
* TERMINAL MAPPING: A = A
*                   B = B
*                   C = C
*                   Y = Y
.SUBCKT AOI21X1_G3 A B C Y 
M19 Y B NET10 0  TSMC20N  L=200E-9 W=2E-6 AD=1E-12 AS=1E-12 PD=5E-6 PS=5E-6 
+M=1 
M20 NET10 A 0 0  TSMC20N  L=200E-9 W=2E-6 AD=1E-12 AS=1E-12 PD=5E-6 PS=5E-6 
+M=1 
M21 Y C 0 0  TSMC20N  L=200E-9 W=1E-6 AD=500E-15 AS=500E-15 PD=3E-6 PS=3E-6 
+M=1 
M16 NET034 A VDD! VDD!  TSMC20P  L=200E-9 W=4E-6 AD=2E-12 AS=2E-12 PD=9E-6 
+PS=9E-6 M=1 
M17 NET034 B VDD! VDD!  TSMC20P  L=200E-9 W=4E-6 AD=2E-12 AS=2E-12 PD=9E-6 
+PS=9E-6 M=1 
M18 Y C NET034 VDD!  TSMC20P  L=200E-9 W=4E-6 AD=2E-12 AS=2E-12 PD=9E-6 
+PS=9E-6 M=1 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS AOI21X1_G3 
* FILE NAME: VITERBI_BMU_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: BMU.
* GENERATED FOR: HSPICES.
* GENERATED ON NOV  7 08:54:36 2007.
   
* TERMINAL MAPPING: BM0<1> = BM0_1
*                   BM0<0> = BM0_0
*                   BM1<1> = BM1_1
*                   BM1<0> = BM1_0
*                   BM2<1> = BM2_1
*                   BM2<0> = BM2_0
*                   BM3<1> = BM3_1
*                   BM3<0> = BM3_0
*                   BM4<1> = BM4_1
*                   BM4<0> = BM4_0
*                   BM5<1> = BM5_1
*                   BM5<0> = BM5_0
*                   BM6<1> = BM6_1
*                   BM6<0> = BM6_0
*                   BM7<1> = BM7_1
*                   BM7<0> = BM7_0
*                   CX0 = CX0
*                   CX1 = CX1
.SUBCKT BMU_G34 BM0_1 BM0_0 BM1_1 BM1_0 BM2_1 BM2_0 BM3_1 BM3_0 BM4_1 BM4_0 
+BM5_1 BM5_0 BM6_1 BM6_0 BM7_1 BM7_0 CX0 CX1 
XU36 CX1 CX0 N2 BM7_0 OAI21X1_G4 
XU38 CX0 CX1 N2 NAND2X1_G9 
XU57 BM3_1 N12 INVX1_G6 
XU58 N12 BM0_1 INVX1_G6 
XU56 N11 BM0_0 INVX1_G6 
XU55 BM3_0 N11 INVX1_G6 
XU53 BM7_1 N10 INVX1_G6 
XU54 N10 BM4_1 INVX1_G6 
XU52 N9 BM4_0 INVX1_G6 
XU51 BM7_0 N9 INVX1_G6 
XU49 BM5_1 N8 INVX1_G6 
XU50 N8 BM6_1 INVX1_G6 
XU48 N7 BM6_0 INVX1_G6 
XU47 BM5_0 N7 INVX1_G6 
XU43 BM3_0 N5 INVX1_G6 
XU44 N5 BM2_0 INVX1_G6 
XU40 N3 BM2_1 INVX1_G6 
XU39 BM1_1 N3 INVX1_G6 
XU45 BM7_0 N6 INVX1_G6 
XU46 N6 BM5_0 INVX1_G6 
XU42 N4 BM1_0 INVX1_G6 
XU37 N2 BM3_1 INVX1_G6 
XU41 BM3_0 N4 INVX1_G6 
XU35 BM7_0 BM3_0 INVX1_G6 
XU33 CX0 N1 INVX1_G6 
XU31 N1 CX1 BM7_1 AND2X1_G8 
XU34 BM3_1 BM3_0 BM1_1 NOR2X1_G7 
XU32 CX1 N1 BM5_1 NOR2X1_G7 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS BMU_G34 
* FILE NAME: VITERBI_SPD_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: SPD.
* GENERATED FOR: HSPICES.
* GENERATED ON NOV  7 08:54:36 2007.
   
* TERMINAL MAPPING: CLK = CLK
*                   D0 = D0
*                   D1 = D1
*                   D2 = D2
*                   D3 = D3
*                   OUT = OUT
*                   PM0<3> = PM0_3
*                   PM0<2> = PM0_2
*                   PM0<1> = PM0_1
*                   PM0<0> = PM0_0
*                   PM1<3> = PM1_3
*                   PM1<2> = PM1_2
*                   PM1<1> = PM1_1
*                   PM1<0> = PM1_0
*                   PM2<3> = PM2_3
*                   PM2<2> = PM2_2
*                   PM2<1> = PM2_1
*                   PM2<0> = PM2_0
*                   PM3<3> = PM3_3
*                   PM3<2> = PM3_2
*                   PM3<1> = PM3_1
*                   PM3<0> = PM3_0
*                   RESET = RESET
.SUBCKT SPD_G33 CLK D0 D1 D2 D3 OUT PM0_3 PM0_2 PM0_1 PM0_0 PM1_3 PM1_2 PM1_1 
+PM1_0 PM2_3 PM2_2 PM2_1 PM2_0 PM3_3 PM3_2 PM3_1 PM3_0 RESET 
XDEMUX1 SELECTORD0 SELECTORD1 SPDU14OUT0 SPDU14OUT1 SPDU14OUT2 SPDU14OUT3 OUT 
+DEMUX_G15 
XSELECTOR1 SELECTORD0 SELECTORD1 PM0_3 PM0_2 PM0_1 PM0_0 PM1_3 PM1_2 PM1_1 
+PM1_0 PM2_3 PM2_2 PM2_1 PM2_0 PM3_3 PM3_2 PM3_1 PM3_0 SELECTOR_G16 
XSPDU13 CLK D0 D1 D2 D3 SPDU12OUT0 SPDU12OUT1 SPDU12OUT2 SPDU12OUT3 SPDU13OUT0 
+SPDU13OUT1 SPDU13OUT2 SPDU13OUT3 RESET SPDU_1_G17 
XSPDU12 CLK D0 D1 D2 D3 SPDU11OUT0 SPDU11OUT1 SPDU11OUT2 SPDU11OUT3 SPDU12OUT0 
+SPDU12OUT1 SPDU12OUT2 SPDU12OUT3 RESET SPDU_2_G18 
XSPDU11 CLK D0 D1 D2 D3 SPDU10OUT0 SPDU10OUT1 SPDU10OUT2 SPDU10OUT3 SPDU11OUT0 
+SPDU11OUT1 SPDU11OUT2 SPDU11OUT3 RESET SPDU_3_G19 
XSPDU10 CLK D0 D1 D2 D3 SPDU9OUT0 SPDU9OUT1 SPDU9OUT2 SPDU9OUT3 SPDU10OUT0 
+SPDU10OUT1 SPDU10OUT2 SPDU10OUT3 RESET SPDU_4_G20 
XSPDU14 CLK D0 D1 D2 D3 SPDU13OUT0 SPDU13OUT1 SPDU13OUT2 SPDU13OUT3 SPDU14OUT0 
+SPDU14OUT1 SPDU14OUT2 SPDU14OUT3 RESET SPDU_0_G21 
XSPDU8 CLK D0 D1 D2 D3 SPDU7OUT0 SPDU7OUT1 SPDU7OUT2 SPDU7OUT3 SPDU8OUT0 
+SPDU8OUT1 SPDU8OUT2 SPDU8OUT3 RESET SPDU_6_G22 
XSPDU7 CLK D0 D1 D2 D3 SPDU6OUT0 SPDU6OUT1 SPDU6OUT2 SPDU6OUT3 SPDU7OUT0 
+SPDU7OUT1 SPDU7OUT2 SPDU7OUT3 RESET SPDU_7_G23 
XSPDU6 CLK D0 D1 D2 D3 SPDU5OUT0 SPDU5OUT1 SPDU5OUT2 SPDU5OUT3 SPDU6OUT0 
+SPDU6OUT1 SPDU6OUT2 SPDU6OUT3 RESET SPDU_8_G24 
XSPDU5 CLK D0 D1 D2 D3 SPDU4OUT0 SPDU4OUT1 SPDU4OUT2 SPDU4OUT3 SPDU5OUT0 
+SPDU5OUT1 SPDU5OUT2 SPDU5OUT3 RESET SPDU_9_G25 
XSPDU9 CLK D0 D1 D2 D3 SPDU8OUT0 SPDU8OUT1 SPDU8OUT2 SPDU8OUT3 SPDU9OUT0 
+SPDU9OUT1 SPDU9OUT2 SPDU9OUT3 RESET SPDU_5_G26 
XSPDU3 CLK D0 D1 D2 D3 SPDU2OUT0 SPDU2OUT1 SPDU2OUT2 SPDU2OUT3 SPDU3OUT0 
+SPDU3OUT1 SPDU3OUT2 SPDU3OUT3 RESET SPDU_11_G27 
XSPDU2 CLK D0 D1 D2 D3 SPDU1OUT0 SPDU1OUT1 SPDU1OUT2 SPDU1OUT3 SPDU2OUT0 
+SPDU2OUT1 SPDU2OUT2 SPDU2OUT3 RESET SPDU_12_G28 
XSPDU1 CLK D0 D1 D2 D3 SPDU0OUT0 SPDU0OUT1 SPDU0OUT2 SPDU0OUT3 SPDU1OUT0 
+SPDU1OUT1 SPDU1OUT2 SPDU1OUT3 RESET SPDU_13_G29 
XSPDU0 CLK D0 D1 D2 D3 GND! GND! VDD! VDD! SPDU0OUT0 SPDU0OUT1 SPDU0OUT2 
+SPDU0OUT3 RESET SPDU_14_G30 
XSPDU4 CLK D0 D1 D2 D3 SPDU3OUT0 SPDU3OUT1 SPDU3OUT2 SPDU3OUT3 SPDU4OUT0 
+SPDU4OUT1 SPDU4OUT2 SPDU4OUT3 RESET SPDU_10_G31 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS SPD_G33 
* FILE NAME: VITERBI_SPDU_10_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: SPDU_10.
* GENERATED FOR: HSPICES.
* GENERATED ON NOV  7 08:54:35 2007.
   
* TERMINAL MAPPING: CLK = CLK
*                   D0 = D0
*                   D1 = D1
*                   D2 = D2
*                   D3 = D3
*                   IN0 = IN0
*                   IN1 = IN1
*                   IN2 = IN2
*                   IN3 = IN3
*                   OUT0 = OUT0
*                   OUT1 = OUT1
*                   OUT2 = OUT2
*                   OUT3 = OUT3
*                   RESET = RESET
.SUBCKT SPDU_10_G31 CLK D0 D1 D2 D3 IN0 IN1 IN2 IN3 OUT0 OUT1 OUT2 OUT3 RESET 
XOUT3_REG CLK OUT3223 OUT3 DFFPOSX1_G14 
XOUT0_REG CLK OUT0205 OUT0 DFFPOSX1_G14 
XOUT2_REG CLK OUT2217 OUT2 DFFPOSX1_G14 
XOUT1_REG CLK OUT1211 OUT1 DFFPOSX1_G14 
XU37 RESET N1 OUT3223 NOR2X1_G7 
XU41 RESET N3 OUT1211 NOR2X1_G7 
XU39 RESET N2 OUT2217 NOR2X1_G7 
XU43 RESET N4 OUT0205 NOR2X1_G7 
XU38 IN3 IN2 D3 N1 MUX2X1_G5 
XU42 IN3 IN2 D1 N3 MUX2X1_G5 
XU44 IN1 IN0 D0 N4 MUX2X1_G5 
XU40 IN1 IN0 D2 N2 MUX2X1_G5 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS SPDU_10_G31 
* FILE NAME: OSU_STDCELLS_OR2X1_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: OR2X1.
* GENERATED FOR: HSPICES.
* GENERATED ON NOV  7 08:54:33 2007.
   
* TERMINAL MAPPING: A = A
*                   B = B
*                   Y = Y
.SUBCKT OR2X1_G13 A B Y 
M14 NET5 B VDD! VDD!  TSMC20P  L=200E-9 W=4E-6 AD=2E-12 AS=2E-12 PD=9E-6 
+PS=9E-6 M=1 
M15 Y NET032 VDD! VDD!  TSMC20P  L=200E-9 W=2E-6 AD=1E-12 AS=1E-12 PD=5E-6 
+PS=5E-6 M=1 
M16 NET032 A NET5 VDD!  TSMC20P  L=200E-9 W=4E-6 AD=2E-12 AS=2E-12 PD=9E-6 
+PS=9E-6 M=1 
M13 NET032 B 0 0  TSMC20N  L=200E-9 W=1E-6 AD=500E-15 AS=500E-15 PD=3E-6 
+PS=3E-6 M=1 
M17 NET032 A 0 0  TSMC20N  L=200E-9 W=1E-6 AD=500E-15 AS=500E-15 PD=3E-6 
+PS=3E-6 M=1 
M18 Y NET032 0 0  TSMC20N  L=200E-9 W=1E-6 AD=500E-15 AS=500E-15 PD=3E-6 
+PS=3E-6 M=1 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS OR2X1_G13 
* FILE NAME: VITERBI_SPDU_3_SCHEMATIC.S.
* SUBCIRCUIT FOR CELL: SPDU_3.
* GENERATED FOR: HSPICES.
* GENERATED ON NOV  7 08:54:34 2007.
   
* TERMINAL MAPPING: CLK = CLK
*                   D0 = D0
*                   D1 = D1
*                   D2 = D2
*                   D3 = D3
*                   IN0 = IN0
*                   IN1 = IN1
*                   IN2 = IN2
*                   IN3 = IN3
*                   OUT0 = OUT0
*                   OUT1 = OUT1
*                   OUT2 = OUT2
*                   OUT3 = OUT3
*                   RESET = RESET
.SUBCKT SPDU_3_G19 CLK D0 D1 D2 D3 IN0 IN1 IN2 IN3 OUT0 OUT1 OUT2 OUT3 RESET 
XOUT0_REG CLK OUT0205 OUT0 DFFPOSX1_G14 
XOUT1_REG CLK OUT1211 OUT1 DFFPOSX1_G14 
XOUT3_REG CLK OUT3223 OUT3 DFFPOSX1_G14 
XOUT2_REG CLK OUT2217 OUT2 DFFPOSX1_G14 
XU41 RESET N3 OUT1211 NOR2X1_G7 
XU39 RESET N2 OUT2217 NOR2X1_G7 
XU43 RESET N4 OUT0205 NOR2X1_G7 
XU37 RESET N1 OUT3223 NOR2X1_G7 
XU38 IN3 IN2 D3 N1 MUX2X1_G5 
XU42 IN3 IN2 D1 N3 MUX2X1_G5 
XU40 IN1 IN0 D2 N2 MUX2X1_G5 
XU44 IN1 IN0 D0 N4 MUX2X1_G5 
   
   
   
* END OF SUBCIRCUIT DEFINITION.
.ENDS SPDU_3_G19 
   
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc20P" PMOS 
.lib "$CDK_DIR/models/hspice/public/publicModel/tsmc20N" NMOS 
   
   
* INCLUDE FILES
   
   
   
   
   
   
* END OF NETLIST
.TEMP    25.0000    
.OP
.save
.OPTION  INGOLD=2 ARTIST=2 PSF=2
+        PROBE=0
.END
