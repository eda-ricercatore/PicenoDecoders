module encoder (b,c);
	output [18:0] c;

	input [7:0] b;

	reg [18:0] c;

	always @(b)
	begin
		c[18] = b[7];
		c[17] = b[6];
		c[16] = b[5];
		c[15] = b[4];
		c[14] = b[3];
		c[13] = b[2];
		c[12] = b[1];
		c[11] = b[0];
		c[10] = b[0] ^ b[2] ^ b[3] ^ b[4] ^ b[5];
		c[9] = b[1] ^ b[4] ^ b[6] ^ b[7];
		c[8] = b[0] ^ b[1] ^ b[3] ^ b[7];
		c[7] = b[0] ^ b[2] ^ b[3];
		c[6] = b[2] ^ b[3] ^ b[5];
		c[5] = b[0] ^ b[1] ^ b[2] ^ b[4] ^ b[7];
		c[4] = b[0] ^ b[1] ^ b[4] ^ b[6];
		c[3] = b[3] ^ b[7];
		c[2] = b[0] ^ b[1] ^ b[3];
		c[1] = b[2] ^ b[3] ^ b[5];
		c[0] = b[1] ^ b[3] ^ b[4] ^ b[5] ^ b[6] ^ b[7];
	end
endmodule
